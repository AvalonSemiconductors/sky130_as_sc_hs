magic
tech sky130A
magscale 1 2
timestamp 1740563454
<< nwell >>
rect -38 262 774 582
<< pwell >>
rect 0 34 736 204
rect 0 22 460 34
rect 26 -20 90 22
<< pmos >>
rect 132 298 162 496
rect 226 298 256 496
rect 356 298 386 496
rect 442 298 472 496
rect 528 298 558 496
rect 614 298 644 496
<< nmoslvt >>
rect 132 48 162 178
rect 226 48 256 178
rect 356 48 386 178
rect 442 48 472 178
rect 528 48 558 178
rect 614 48 644 178
<< ndiff >>
rect 74 164 132 178
rect 74 130 87 164
rect 121 130 132 164
rect 74 48 132 130
rect 162 48 226 178
rect 256 94 356 178
rect 256 60 311 94
rect 345 60 356 94
rect 256 48 356 60
rect 386 170 442 178
rect 386 136 397 170
rect 431 136 442 170
rect 386 48 442 136
rect 472 166 528 178
rect 472 60 483 166
rect 517 60 528 166
rect 472 48 528 60
rect 558 170 614 178
rect 558 136 569 170
rect 603 136 614 170
rect 558 48 614 136
rect 644 170 709 178
rect 644 56 660 170
rect 694 56 709 170
rect 644 48 709 56
<< pdiff >>
rect 72 488 132 496
rect 72 316 85 488
rect 119 316 132 488
rect 72 298 132 316
rect 162 434 226 496
rect 162 328 176 434
rect 210 328 226 434
rect 162 298 226 328
rect 256 488 356 496
rect 256 420 286 488
rect 320 420 356 488
rect 256 298 356 420
rect 386 476 442 496
rect 386 306 397 476
rect 431 306 442 476
rect 386 298 442 306
rect 472 484 528 496
rect 472 338 483 484
rect 517 338 528 484
rect 472 298 528 338
rect 558 476 614 496
rect 558 306 569 476
rect 603 306 614 476
rect 558 298 614 306
rect 644 488 709 496
rect 644 308 656 488
rect 690 308 709 488
rect 644 298 709 308
<< ndiffc >>
rect 87 130 121 164
rect 311 60 345 94
rect 397 136 431 170
rect 483 60 517 166
rect 569 136 603 170
rect 660 56 694 170
<< pdiffc >>
rect 85 316 119 488
rect 176 328 210 434
rect 286 420 320 488
rect 397 306 431 476
rect 483 338 517 484
rect 569 306 603 476
rect 656 308 690 488
<< poly >>
rect 132 496 162 522
rect 226 496 256 522
rect 356 496 386 522
rect 442 496 472 522
rect 528 496 558 522
rect 614 496 644 522
rect 132 266 162 298
rect 226 266 256 298
rect 356 266 386 298
rect 116 250 170 266
rect 116 216 126 250
rect 160 216 170 250
rect 116 198 170 216
rect 222 250 276 266
rect 222 216 232 250
rect 266 216 276 250
rect 222 198 276 216
rect 318 264 386 266
rect 442 264 472 298
rect 318 258 472 264
rect 528 258 558 298
rect 318 250 558 258
rect 318 216 328 250
rect 362 234 558 250
rect 614 234 644 298
rect 362 222 644 234
rect 362 216 472 222
rect 318 198 472 216
rect 132 178 162 198
rect 226 178 256 198
rect 356 178 386 198
rect 442 178 472 198
rect 528 198 644 222
rect 528 178 558 198
rect 614 178 644 198
rect 132 22 162 48
rect 226 22 256 48
rect 356 22 386 48
rect 442 22 472 48
rect 528 22 558 48
rect 614 22 644 48
<< polycont >>
rect 126 216 160 250
rect 232 216 266 250
rect 328 216 362 250
<< locali >>
rect 0 561 736 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 526 736 527
rect 85 488 119 526
rect 286 488 320 526
rect 85 300 119 316
rect 176 434 210 450
rect 286 402 320 420
rect 397 476 431 492
rect 210 328 362 346
rect 176 312 362 328
rect 68 250 170 266
rect 68 216 126 250
rect 160 216 170 250
rect 68 198 170 216
rect 222 250 276 278
rect 222 216 232 250
rect 266 216 276 250
rect 222 198 276 216
rect 328 250 362 312
rect 328 164 362 216
rect 71 130 87 164
rect 121 130 362 164
rect 483 484 517 526
rect 483 322 517 338
rect 569 476 603 492
rect 397 296 431 306
rect 397 270 460 296
rect 569 270 603 306
rect 656 488 690 526
rect 656 292 690 308
rect 397 234 603 270
rect 397 214 460 234
rect 397 170 431 214
rect 397 120 431 136
rect 483 166 517 182
rect 294 94 362 96
rect 294 60 311 94
rect 345 60 362 94
rect 569 170 603 234
rect 569 120 603 136
rect 660 170 694 186
rect 311 21 345 60
rect 483 21 517 60
rect 660 21 694 56
rect 0 17 736 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 68 221 102 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 85 238 85 238 0 FreeSans 200 0 0 0 A
flabel locali s 238 221 272 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 255 238 255 238 0 FreeSans 200 0 0 0 B
flabel locali s 408 221 442 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 425 238 425 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__and2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 736 220
string MASKHINTS_NSDM 0 -38 736 209
string MASKHINTS_PSDM 0 273 736 582
<< end >>
