.option method=key
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt_mm
.option wnflag=1

.include ./sky130_as_sc_hs__nand2_1.spice

VDD VPWR 0 1.8V
VSS VGND 0 0V

R111 VNB GND 0
R112 VPB VPWR 0
R113 GND VGND 0

Va A GND PULSE( 0 1.8 0 0.1ns 0.1ns 5ns 10ns )
Vb B GND PULSE( 0 1.8 0 0.1ns 0.1ns 10ns 20ns )

.tran 1n 50n

.control
run
plot v(A)+2 v(B) v(Y)
.endc
.end
