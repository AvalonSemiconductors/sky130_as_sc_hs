magic
tech sky130A
magscale 1 2
timestamp 1733756788
<< nwell >>
rect -38 262 314 582
<< pwell >>
rect 2 44 274 204
rect 26 -15 76 44
rect 26 -20 66 -15
<< poly >>
rect 60 478 208 494
rect 60 384 156 478
rect 198 384 208 478
rect 60 346 208 384
rect 60 304 208 336
rect 60 92 72 304
rect 196 92 208 304
rect 60 48 208 92
<< polycont >>
rect 156 384 198 478
rect 72 92 196 304
<< rmp >>
rect 60 336 208 346
<< locali >>
rect 0 561 276 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 526 276 527
rect 146 478 208 526
rect 146 384 156 478
rect 198 384 208 478
rect 146 368 208 384
rect 60 304 208 326
rect 60 92 72 304
rect 196 92 208 304
rect 60 76 208 92
rect 0 17 276 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel comment s 0 0 0 0 4 tieh
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 276 48 1 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 153 272 187 306 0 FreeSans 200 0 0 0 ONE
port 5 nsew signal output
flabel locali s 170 289 170 289 0 FreeSans 200 0 0 0 ONE
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__tieh.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 276 227
string MASKHINTS_NSDM 0 -38 276 203
string MASKHINTS_PSDM 0 272 276 582
<< end >>
