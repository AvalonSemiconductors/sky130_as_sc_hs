magic
tech sky130A
magscale 1 2
timestamp 1740335508
<< nwell >>
rect -38 262 866 582
<< pwell >>
rect 0 26 828 204
rect 22 24 90 26
rect 22 22 110 24
rect 168 22 198 24
rect 256 22 286 24
rect 344 22 374 24
rect 432 22 462 24
rect 519 22 549 24
rect 605 22 635 24
rect 691 22 721 24
rect 22 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 168 298 198 496
rect 256 298 286 496
rect 344 298 374 496
rect 432 298 462 496
rect 519 298 549 496
rect 605 298 635 496
rect 691 298 721 496
<< nmoslvt >>
rect 80 48 110 178
rect 168 48 198 178
rect 256 48 286 178
rect 344 48 374 178
rect 432 48 462 178
rect 519 48 549 178
rect 605 48 635 178
rect 691 48 721 178
<< ndiff >>
rect 27 140 80 178
rect 27 76 35 140
rect 69 76 80 140
rect 27 48 80 76
rect 110 170 168 178
rect 110 72 121 170
rect 155 72 168 170
rect 110 48 168 72
rect 198 150 256 178
rect 198 58 209 150
rect 243 58 256 150
rect 198 48 256 58
rect 286 150 344 178
rect 286 116 298 150
rect 332 116 344 150
rect 286 48 344 116
rect 374 106 432 178
rect 374 72 386 106
rect 420 72 432 106
rect 374 48 432 72
rect 462 164 519 178
rect 462 130 474 164
rect 508 130 519 164
rect 462 48 519 130
rect 549 166 605 178
rect 549 57 560 166
rect 594 57 605 166
rect 549 48 605 57
rect 635 152 691 178
rect 635 118 646 152
rect 680 118 691 152
rect 635 48 691 118
rect 721 170 801 178
rect 721 57 736 170
rect 770 57 801 170
rect 721 48 801 57
<< pdiff >>
rect 27 484 80 496
rect 27 350 35 484
rect 69 350 80 484
rect 27 298 80 350
rect 110 476 168 496
rect 110 331 121 476
rect 155 331 168 476
rect 110 298 168 331
rect 198 488 256 496
rect 198 346 209 488
rect 243 346 256 488
rect 198 298 256 346
rect 286 476 344 496
rect 286 354 298 476
rect 332 354 344 476
rect 286 298 344 354
rect 374 474 432 496
rect 374 406 386 474
rect 420 406 432 474
rect 374 298 432 406
rect 462 474 519 496
rect 462 354 474 474
rect 508 354 519 474
rect 462 298 519 354
rect 549 488 605 496
rect 549 342 560 488
rect 594 342 605 488
rect 549 298 605 342
rect 635 474 691 496
rect 635 331 646 474
rect 680 331 691 474
rect 635 298 691 331
rect 721 488 801 496
rect 721 342 734 488
rect 768 342 801 488
rect 721 298 801 342
<< ndiffc >>
rect 35 76 69 140
rect 121 72 155 170
rect 209 58 243 150
rect 298 116 332 150
rect 386 72 420 106
rect 474 130 508 164
rect 560 57 594 166
rect 646 118 680 152
rect 736 57 770 170
<< pdiffc >>
rect 35 350 69 484
rect 121 331 155 476
rect 209 346 243 488
rect 298 354 332 476
rect 386 406 420 474
rect 474 354 508 474
rect 560 342 594 488
rect 646 331 680 474
rect 734 342 768 488
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 519 496 549 522
rect 605 496 635 522
rect 691 496 721 522
rect 80 282 110 298
rect 168 282 198 298
rect 80 266 198 282
rect 256 280 286 298
rect 344 280 374 298
rect 432 280 462 298
rect 519 280 549 298
rect 256 270 549 280
rect 40 250 198 266
rect 40 216 50 250
rect 84 226 198 250
rect 84 216 110 226
rect 40 200 110 216
rect 80 178 110 200
rect 168 178 198 226
rect 240 260 549 270
rect 605 262 635 298
rect 691 262 721 298
rect 605 260 721 262
rect 240 250 721 260
rect 240 216 250 250
rect 284 230 721 250
rect 284 216 296 230
rect 240 204 296 216
rect 240 200 286 204
rect 256 178 286 200
rect 344 178 374 230
rect 432 178 462 230
rect 519 178 549 230
rect 605 178 635 230
rect 691 178 721 230
rect 80 22 110 48
rect 168 22 198 48
rect 256 22 286 48
rect 344 22 374 48
rect 432 22 462 48
rect 519 22 549 48
rect 605 22 635 48
rect 691 22 721 48
<< polycont >>
rect 50 216 84 250
rect 250 216 284 250
<< locali >>
rect 0 561 828 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 526 828 527
rect 35 484 69 526
rect 35 334 69 350
rect 120 476 156 492
rect 120 331 121 476
rect 155 331 156 476
rect 31 250 84 296
rect 31 216 50 250
rect 31 192 84 216
rect 120 284 156 331
rect 209 488 243 526
rect 209 330 243 346
rect 298 476 332 492
rect 386 474 420 526
rect 386 390 420 406
rect 474 474 508 490
rect 332 354 356 372
rect 298 338 356 354
rect 322 292 356 338
rect 474 292 508 354
rect 560 488 594 526
rect 560 326 594 342
rect 646 474 680 490
rect 646 292 680 331
rect 734 488 768 526
rect 734 326 768 342
rect 120 250 284 284
rect 120 244 250 250
rect 120 170 156 244
rect 238 216 250 244
rect 238 200 284 216
rect 322 252 680 292
rect 322 188 356 252
rect 35 140 69 158
rect 35 21 69 76
rect 120 72 121 170
rect 155 72 156 170
rect 318 166 356 188
rect 120 56 156 72
rect 209 150 243 166
rect 298 154 356 166
rect 474 238 680 252
rect 474 164 508 238
rect 298 150 352 154
rect 332 130 352 150
rect 298 100 332 116
rect 386 106 420 122
rect 474 114 508 130
rect 560 166 594 182
rect 209 21 243 58
rect 386 21 420 72
rect 646 152 680 238
rect 646 102 680 118
rect 736 170 770 190
rect 560 21 594 57
rect 736 21 770 57
rect 0 17 828 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_6
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali 357 255 391 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 374 272 374 272 0 FreeSans 200 0 0 0 Y
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_6.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 828 216
string MASKHINTS_NSDM 0 -38 828 204
string MASKHINTS_PSDM 0 272 828 582
<< end >>
