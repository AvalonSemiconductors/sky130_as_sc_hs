magic
tech sky130A
magscale 1 2
timestamp 1736644844
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 0 -4 460 204
rect 26 -20 90 -4
<< pmos >>
rect 80 314 110 496
rect 166 314 196 496
rect 252 314 282 496
rect 338 314 368 496
<< nmoslvt >>
rect 80 49 110 176
rect 166 49 196 176
rect 252 49 282 176
rect 338 49 368 176
<< ndiff >>
rect 27 156 80 176
rect 27 64 35 156
rect 69 64 80 156
rect 27 49 80 64
rect 110 154 166 176
rect 110 76 121 154
rect 155 76 166 154
rect 110 49 166 76
rect 196 92 252 176
rect 196 58 207 92
rect 241 58 252 92
rect 196 49 252 58
rect 282 150 338 176
rect 282 72 293 150
rect 327 72 338 150
rect 282 49 338 72
rect 368 92 433 176
rect 368 58 380 92
rect 414 58 433 92
rect 368 49 433 58
<< pdiff >>
rect 27 476 80 496
rect 27 344 35 476
rect 69 344 80 476
rect 27 314 80 344
rect 110 486 166 496
rect 110 410 121 486
rect 155 410 166 486
rect 110 314 166 410
rect 196 476 252 496
rect 196 340 207 476
rect 241 340 252 476
rect 196 314 252 340
rect 282 398 338 496
rect 282 322 293 398
rect 327 322 338 398
rect 282 314 338 322
rect 368 476 433 496
rect 368 400 386 476
rect 420 400 433 476
rect 368 314 433 400
<< ndiffc >>
rect 35 64 69 156
rect 121 76 155 154
rect 207 58 241 92
rect 293 72 327 150
rect 380 58 414 92
<< pdiffc >>
rect 35 344 69 476
rect 121 410 155 486
rect 207 340 241 476
rect 293 322 327 398
rect 386 400 420 476
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 80 268 110 314
rect 166 268 196 314
rect 252 268 282 314
rect 338 268 368 314
rect 62 250 196 268
rect 62 216 78 250
rect 180 216 196 250
rect 62 200 196 216
rect 238 252 370 268
rect 238 218 254 252
rect 306 218 370 252
rect 238 200 370 218
rect 80 176 110 200
rect 166 176 196 200
rect 252 176 282 200
rect 338 176 368 200
rect 80 23 110 49
rect 166 23 196 49
rect 252 23 282 49
rect 338 23 368 49
<< polycont >>
rect 78 216 180 250
rect 254 218 306 252
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 30 476 76 492
rect 30 344 35 476
rect 69 360 76 476
rect 110 486 166 526
rect 110 410 121 486
rect 155 410 166 486
rect 110 394 166 410
rect 200 476 432 492
rect 200 360 207 476
rect 69 344 207 360
rect 30 340 207 344
rect 241 448 386 476
rect 241 340 248 448
rect 30 314 248 340
rect 284 398 336 414
rect 284 322 293 398
rect 327 350 336 398
rect 382 400 386 448
rect 420 400 432 476
rect 382 384 432 400
rect 327 322 432 350
rect 284 304 432 322
rect 62 250 196 268
rect 62 216 78 250
rect 180 216 196 250
rect 62 212 196 216
rect 238 252 322 268
rect 238 218 254 252
rect 306 218 322 252
rect 238 212 322 218
rect 356 178 432 304
rect 35 156 69 172
rect 35 21 69 64
rect 114 154 432 178
rect 114 76 121 154
rect 155 150 432 154
rect 155 142 293 150
rect 155 76 158 142
rect 114 56 158 76
rect 207 92 241 108
rect 207 21 241 58
rect 288 72 293 142
rect 327 142 432 150
rect 327 72 332 142
rect 288 56 332 72
rect 380 92 414 108
rect 380 21 414 58
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 A
flabel locali 255 221 289 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 272 238 272 238 0 FreeSans 200 0 0 0 B
flabel locali 391 187 425 221 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 408 204 408 204 0 FreeSans 200 0 0 0 Y
flabel locali 391 289 425 323 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 408 306 408 306 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 214
string MASKHINTS_NSDM 0 -38 460 201
string MASKHINTS_PSDM 0 289 460 582
<< end >>
