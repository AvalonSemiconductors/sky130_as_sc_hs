magic
tech sky130A
magscale 1 2
timestamp 1740391790
<< nwell >>
rect -38 262 1234 582
<< pwell >>
rect 0 26 1196 204
rect 0 24 920 26
rect 930 24 1196 26
rect 0 22 736 24
rect 782 22 812 24
rect 904 22 934 24
rect 990 22 1020 24
rect 1076 22 1106 24
rect 26 -20 90 22
<< pmos >>
rect 80 347 110 496
rect 166 347 196 496
rect 284 298 314 496
rect 434 298 464 496
rect 672 298 702 496
rect 782 298 812 496
rect 904 298 934 496
rect 990 298 1020 496
rect 1076 298 1106 496
<< nmoslvt >>
rect 80 48 110 166
rect 176 48 206 166
rect 284 48 314 178
rect 544 48 574 178
rect 672 48 702 178
rect 782 48 812 178
rect 904 48 934 178
rect 990 48 1020 178
rect 1076 48 1106 178
<< ndiff >>
rect 230 166 284 178
rect 27 154 80 166
rect 27 72 35 154
rect 69 72 80 154
rect 27 48 80 72
rect 110 102 176 166
rect 110 68 121 102
rect 155 68 176 102
rect 110 48 176 68
rect 206 48 284 166
rect 314 150 544 178
rect 314 116 329 150
rect 363 116 544 150
rect 314 90 544 116
rect 314 56 386 90
rect 420 56 544 90
rect 314 48 544 56
rect 574 148 672 178
rect 574 114 624 148
rect 658 114 672 148
rect 574 48 672 114
rect 702 150 782 178
rect 702 58 718 150
rect 752 58 782 150
rect 702 48 782 58
rect 812 166 904 178
rect 812 132 858 166
rect 892 132 904 166
rect 812 48 904 132
rect 934 164 990 178
rect 934 58 945 164
rect 979 58 990 164
rect 934 48 990 58
rect 1020 170 1076 178
rect 1020 136 1031 170
rect 1065 136 1076 170
rect 1020 48 1076 136
rect 1106 164 1160 178
rect 1106 62 1117 164
rect 1151 62 1160 164
rect 1106 48 1160 62
<< pdiff >>
rect 27 472 80 496
rect 27 438 35 472
rect 69 438 80 472
rect 27 347 80 438
rect 110 474 166 496
rect 110 440 121 474
rect 155 440 166 474
rect 110 347 166 440
rect 196 347 284 496
rect 230 298 284 347
rect 314 446 434 496
rect 314 412 356 446
rect 390 412 434 446
rect 314 298 434 412
rect 464 346 672 496
rect 464 312 488 346
rect 522 312 564 346
rect 598 312 672 346
rect 464 298 672 312
rect 702 488 782 496
rect 702 454 716 488
rect 750 454 782 488
rect 702 298 782 454
rect 812 470 904 496
rect 812 322 858 470
rect 892 322 904 470
rect 812 298 904 322
rect 934 488 990 496
rect 934 320 945 488
rect 979 320 990 488
rect 934 298 990 320
rect 1020 474 1076 496
rect 1020 306 1031 474
rect 1065 306 1076 474
rect 1020 298 1076 306
rect 1106 484 1160 496
rect 1106 312 1117 484
rect 1151 312 1160 484
rect 1106 298 1160 312
<< ndiffc >>
rect 35 72 69 154
rect 121 68 155 102
rect 329 116 363 150
rect 386 56 420 90
rect 624 114 658 148
rect 718 58 752 150
rect 858 132 892 166
rect 945 58 979 164
rect 1031 136 1065 170
rect 1117 62 1151 164
<< pdiffc >>
rect 35 438 69 472
rect 121 440 155 474
rect 356 412 390 446
rect 488 312 522 346
rect 564 312 598 346
rect 716 454 750 488
rect 858 322 892 470
rect 945 320 979 488
rect 1031 306 1065 474
rect 1117 312 1151 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 284 496 314 522
rect 434 496 464 522
rect 672 496 702 522
rect 782 496 812 522
rect 904 496 934 522
rect 990 496 1020 522
rect 1076 496 1106 522
rect 80 332 110 347
rect 166 332 196 347
rect 80 302 196 332
rect 80 296 133 302
rect 79 280 133 296
rect 79 246 89 280
rect 123 246 133 280
rect 284 266 314 298
rect 79 230 133 246
rect 176 250 242 260
rect 80 166 110 230
rect 176 216 192 250
rect 226 216 242 250
rect 176 206 242 216
rect 284 250 392 266
rect 284 216 346 250
rect 380 216 392 250
rect 176 166 206 206
rect 284 200 392 216
rect 434 260 464 298
rect 672 266 702 298
rect 782 266 812 298
rect 904 266 934 298
rect 990 266 1020 298
rect 1076 266 1106 298
rect 434 250 502 260
rect 434 216 450 250
rect 484 216 502 250
rect 434 206 502 216
rect 544 250 598 266
rect 544 216 554 250
rect 588 216 598 250
rect 544 200 598 216
rect 672 250 740 266
rect 672 216 692 250
rect 726 216 740 250
rect 672 200 740 216
rect 782 250 1106 266
rect 782 216 792 250
rect 826 216 1106 250
rect 782 200 1106 216
rect 284 178 314 200
rect 544 178 574 200
rect 672 178 702 200
rect 782 178 812 200
rect 904 178 934 200
rect 990 178 1020 200
rect 1076 178 1106 200
rect 80 22 110 48
rect 176 22 206 48
rect 284 22 314 48
rect 544 22 574 48
rect 672 22 702 48
rect 782 22 812 48
rect 904 22 934 48
rect 990 22 1020 48
rect 1076 22 1106 48
<< polycont >>
rect 89 246 123 280
rect 192 216 226 250
rect 346 216 380 250
rect 450 216 484 250
rect 554 216 588 250
rect 692 216 726 250
rect 792 216 826 250
<< locali >>
rect 0 561 1196 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 526 1196 527
rect 20 472 69 488
rect 20 418 35 472
rect 20 404 69 418
rect 121 474 155 526
rect 716 488 750 526
rect 945 488 979 526
rect 121 412 155 440
rect 278 412 356 446
rect 390 412 682 446
rect 716 438 750 454
rect 858 470 894 486
rect 20 186 55 404
rect 89 336 210 370
rect 89 280 136 336
rect 123 246 136 280
rect 89 220 136 246
rect 176 250 242 252
rect 176 216 192 250
rect 226 216 242 250
rect 176 208 242 216
rect 176 186 210 208
rect 20 154 210 186
rect 20 150 35 154
rect 69 152 210 154
rect 278 166 312 412
rect 648 402 682 412
rect 648 368 808 402
rect 472 334 488 346
rect 358 312 488 334
rect 522 312 564 346
rect 598 334 616 346
rect 598 312 658 334
rect 358 300 658 312
rect 358 266 392 300
rect 346 250 392 266
rect 380 216 392 250
rect 346 200 392 216
rect 434 250 502 260
rect 484 216 502 250
rect 434 214 502 216
rect 544 250 590 266
rect 544 216 554 250
rect 588 216 590 250
rect 544 200 590 216
rect 544 180 578 200
rect 426 166 578 180
rect 278 150 363 166
rect 278 128 329 150
rect 35 56 69 72
rect 121 102 155 118
rect 121 21 155 68
rect 460 146 578 166
rect 624 148 658 300
rect 774 266 808 368
rect 892 322 894 470
rect 858 306 894 322
rect 860 268 908 306
rect 945 304 979 320
rect 1031 474 1065 490
rect 1031 268 1065 306
rect 1117 484 1151 526
rect 1117 296 1151 312
rect 692 250 740 266
rect 726 216 740 250
rect 692 200 740 216
rect 774 250 826 266
rect 774 216 792 250
rect 774 200 826 216
rect 860 226 1065 268
rect 860 182 908 226
rect 858 166 894 182
rect 329 90 363 116
rect 624 98 658 114
rect 718 150 752 166
rect 329 56 386 90
rect 420 56 436 90
rect 892 132 894 166
rect 858 116 894 132
rect 945 164 979 180
rect 718 21 752 58
rect 1031 170 1065 226
rect 1031 120 1065 136
rect 1117 164 1151 180
rect 945 21 979 58
rect 1117 21 1151 62
rect 0 17 1196 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 35 438 69 452
rect 35 418 69 438
rect 210 336 244 370
rect 434 216 450 250
rect 450 216 468 250
rect 426 132 460 166
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 22 454 80 458
rect 22 452 466 454
rect 22 418 35 452
rect 69 418 466 452
rect 22 416 466 418
rect 22 412 80 416
rect 198 370 282 382
rect 198 336 210 370
rect 244 336 282 370
rect 198 328 282 336
rect 248 182 282 328
rect 434 256 466 416
rect 422 250 480 256
rect 422 216 434 250
rect 468 216 480 250
rect 422 210 480 216
rect 248 166 472 182
rect 248 146 426 166
rect 414 132 426 146
rect 460 132 472 166
rect 414 126 472 132
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 102 238 136 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 697 221 731 255 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel locali 714 238 714 238 0 FreeSans 200 0 0 0 B
flabel locali 867 221 901 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 884 238 884 238 0 FreeSans 200 0 0 0 Y
flabel polycont 119 255 119 255 0 FreeSans 200 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__xnor2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1196 214
string MASKHINTS_NSDM 0 -38 1196 204
string MASKHINTS_PSDM 0 272 1196 582
<< end >>
