magic
tech sky130A
magscale 1 2
timestamp 1733931690
<< nwell >>
rect -38 262 1052 582
<< pwell >>
rect 20 44 1012 204
rect 20 -15 82 44
rect 20 -20 74 -15
<< pmos >>
rect 81 298 111 496
rect 168 298 198 496
rect 256 298 286 496
rect 344 298 374 496
rect 432 298 462 496
rect 524 298 554 496
rect 612 298 642 496
rect 700 298 730 496
rect 788 298 818 496
rect 876 298 906 496
<< nmoslvt >>
rect 81 47 111 134
rect 168 47 198 134
rect 256 47 286 134
rect 344 47 374 134
rect 432 47 462 134
rect 524 47 554 134
rect 612 47 642 134
rect 700 47 730 134
rect 788 47 818 134
rect 876 47 906 134
<< ndiff >>
rect 28 116 81 134
rect 28 64 36 116
rect 70 64 81 116
rect 28 47 81 64
rect 111 126 168 134
rect 111 72 122 126
rect 156 72 168 126
rect 111 47 168 72
rect 198 94 256 134
rect 198 56 210 94
rect 244 56 256 94
rect 198 47 256 56
rect 286 126 344 134
rect 286 72 298 126
rect 332 72 344 126
rect 286 47 344 72
rect 374 94 432 134
rect 374 56 386 94
rect 420 56 432 94
rect 374 47 432 56
rect 462 126 524 134
rect 462 72 478 126
rect 512 72 524 126
rect 462 47 524 72
rect 554 96 612 134
rect 554 56 566 96
rect 600 56 612 96
rect 554 47 612 56
rect 642 126 700 134
rect 642 72 654 126
rect 688 72 700 126
rect 642 47 700 72
rect 730 96 788 134
rect 730 56 742 96
rect 776 56 788 96
rect 730 47 788 56
rect 818 126 876 134
rect 818 72 830 126
rect 864 72 876 126
rect 818 47 876 72
rect 906 96 964 134
rect 906 56 918 96
rect 952 56 964 96
rect 906 47 964 56
<< pdiff >>
rect 28 480 81 496
rect 28 324 36 480
rect 70 324 81 480
rect 28 298 81 324
rect 111 476 168 496
rect 111 334 122 476
rect 156 334 168 476
rect 111 298 168 334
rect 198 482 256 496
rect 198 386 210 482
rect 244 386 256 482
rect 198 298 256 386
rect 286 476 344 496
rect 286 336 298 476
rect 332 336 344 476
rect 286 298 344 336
rect 374 484 432 496
rect 374 386 386 484
rect 420 386 432 484
rect 374 298 432 386
rect 462 476 524 496
rect 462 334 478 476
rect 512 334 524 476
rect 462 298 524 334
rect 554 484 612 496
rect 554 386 566 484
rect 600 386 612 484
rect 554 298 612 386
rect 642 476 700 496
rect 642 334 654 476
rect 688 334 700 476
rect 642 298 700 334
rect 730 484 788 496
rect 730 386 742 484
rect 776 386 788 484
rect 730 298 788 386
rect 818 476 876 496
rect 818 334 830 476
rect 864 334 876 476
rect 818 298 876 334
rect 906 484 960 496
rect 906 386 918 484
rect 952 386 960 484
rect 906 298 960 386
<< ndiffc >>
rect 36 64 70 116
rect 122 72 156 126
rect 210 56 244 94
rect 298 72 332 126
rect 386 56 420 94
rect 478 72 512 126
rect 566 56 600 96
rect 654 72 688 126
rect 742 56 776 96
rect 830 72 864 126
rect 918 56 952 96
<< pdiffc >>
rect 36 324 70 480
rect 122 334 156 476
rect 210 386 244 482
rect 298 336 332 476
rect 386 386 420 484
rect 478 334 512 476
rect 566 386 600 484
rect 654 334 688 476
rect 742 386 776 484
rect 830 334 864 476
rect 918 386 952 484
<< poly >>
rect 81 496 111 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 524 496 554 522
rect 612 496 642 522
rect 700 496 730 522
rect 788 496 818 522
rect 876 496 906 522
rect 81 268 111 298
rect 168 268 198 298
rect 60 248 198 268
rect 60 214 76 248
rect 180 214 198 248
rect 60 204 198 214
rect 81 134 111 204
rect 168 134 198 204
rect 256 262 286 298
rect 344 262 374 298
rect 432 262 462 298
rect 524 262 554 298
rect 612 262 642 298
rect 700 262 730 298
rect 788 262 818 298
rect 876 262 906 298
rect 256 248 906 262
rect 256 214 272 248
rect 760 214 906 248
rect 256 204 906 214
rect 256 134 286 204
rect 344 134 374 204
rect 432 134 462 204
rect 524 134 554 204
rect 612 134 642 204
rect 700 134 730 204
rect 788 134 818 204
rect 876 134 906 204
rect 81 21 111 47
rect 168 21 198 47
rect 256 21 286 47
rect 344 21 374 47
rect 432 21 462 47
rect 524 21 554 47
rect 612 21 642 47
rect 700 21 730 47
rect 788 21 818 47
rect 876 21 906 47
<< polycont >>
rect 76 214 180 248
rect 272 214 760 248
<< locali >>
rect 0 561 1014 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1014 561
rect 0 526 1014 527
rect 26 480 80 526
rect 26 324 36 480
rect 70 324 80 480
rect 26 308 80 324
rect 114 476 164 492
rect 114 334 122 476
rect 156 336 164 476
rect 200 482 254 526
rect 200 386 210 482
rect 244 386 254 482
rect 200 370 254 386
rect 298 476 342 492
rect 332 336 342 476
rect 376 484 430 526
rect 376 386 386 484
rect 420 386 430 484
rect 376 370 430 386
rect 478 476 522 492
rect 156 334 264 336
rect 114 302 264 334
rect 298 334 478 336
rect 512 336 522 476
rect 556 484 610 526
rect 556 386 566 484
rect 600 386 610 484
rect 556 370 610 386
rect 644 476 698 492
rect 644 336 654 476
rect 512 334 654 336
rect 688 336 698 476
rect 732 484 786 526
rect 732 386 742 484
rect 776 386 786 484
rect 732 370 786 386
rect 820 476 874 492
rect 820 336 830 476
rect 688 334 830 336
rect 864 336 874 476
rect 908 484 962 526
rect 908 386 918 484
rect 952 386 962 484
rect 908 370 962 386
rect 864 334 984 336
rect 298 302 984 334
rect 230 268 264 302
rect 26 248 196 268
rect 26 214 76 248
rect 180 214 196 248
rect 230 248 776 268
rect 230 214 272 248
rect 760 214 776 248
rect 26 168 80 214
rect 230 180 264 214
rect 810 180 984 302
rect 114 146 264 180
rect 298 146 984 180
rect 28 116 78 134
rect 28 64 36 116
rect 70 64 78 116
rect 28 21 78 64
rect 114 126 164 146
rect 114 72 122 126
rect 156 72 164 126
rect 298 126 340 146
rect 114 56 164 72
rect 202 94 252 110
rect 202 56 210 94
rect 244 56 252 94
rect 332 72 340 126
rect 478 126 520 146
rect 298 56 340 72
rect 378 94 428 110
rect 378 56 386 94
rect 420 56 428 94
rect 512 72 520 126
rect 646 126 696 146
rect 478 56 520 72
rect 558 96 608 112
rect 558 56 566 96
rect 600 56 608 96
rect 646 72 654 126
rect 688 72 696 126
rect 822 126 872 146
rect 646 56 696 72
rect 734 96 784 112
rect 734 56 742 96
rect 776 56 784 96
rect 822 72 830 126
rect 864 72 872 126
rect 822 56 872 72
rect 910 96 960 112
rect 910 56 918 96
rect 952 56 960 96
rect 202 21 252 56
rect 378 21 428 56
rect 558 21 608 56
rect 734 21 784 56
rect 910 21 960 56
rect 0 17 1012 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1014 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1014 561
rect 0 496 1014 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel comment s 0 0 0 0 4 clkbuff_8
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 0 496 1014 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali 935 187 969 221 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel locali 952 204 952 204 0 FreeSans 200 0 0 0 Y
flabel locali 816 187 850 221 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel locali 833 204 833 204 0 FreeSans 200 0 0 0 Y
flabel locali 816 289 850 323 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel locali 833 306 833 306 0 FreeSans 200 0 0 0 Y
flabel locali 935 289 969 323 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel locali 952 306 952 306 0 FreeSans 200 0 0 0 Y
flabel locali 34 170 68 204 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 51 187 51 187 0 FreeSans 200 0 0 0 A
flabel locali 102 221 136 255 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 119 238 119 238 0 FreeSans 200 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__clkbuff_8.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
