magic
tech sky130A
magscale 1 2
timestamp 1733959029
<< nwell >>
rect -38 262 1510 582
<< pwell >>
rect 20 44 1424 204
rect 20 -15 82 44
rect 20 -20 74 -15
<< nmos >>
rect 81 50 111 158
rect 168 50 198 158
rect 256 50 286 158
rect 344 50 374 158
rect 432 50 462 158
rect 524 50 554 158
rect 612 50 642 158
rect 700 50 730 158
rect 788 50 818 158
rect 876 50 906 158
rect 964 50 994 158
rect 1052 50 1082 158
rect 1140 50 1170 158
rect 1230 50 1260 158
rect 1318 50 1348 158
<< pmos >>
rect 81 352 111 496
rect 168 352 198 496
rect 256 352 286 496
rect 344 352 374 496
rect 432 352 462 496
rect 524 352 554 496
rect 612 352 642 496
rect 700 352 730 496
rect 788 352 818 496
rect 876 352 906 496
rect 964 352 994 496
rect 1052 352 1082 496
rect 1140 352 1170 496
rect 1230 352 1260 496
rect 1318 352 1348 496
<< ndiff >>
rect 28 132 81 158
rect 28 64 36 132
rect 70 64 81 132
rect 28 50 81 64
rect 111 150 168 158
rect 111 72 122 150
rect 156 72 168 150
rect 111 50 168 72
rect 198 124 256 158
rect 198 64 210 124
rect 244 64 256 124
rect 198 50 256 64
rect 286 150 344 158
rect 286 72 298 150
rect 332 72 344 150
rect 286 50 344 72
rect 374 124 432 158
rect 374 64 386 124
rect 420 64 432 124
rect 374 50 432 64
rect 462 150 524 158
rect 462 72 478 150
rect 512 72 524 150
rect 462 50 524 72
rect 554 124 612 158
rect 554 64 566 124
rect 600 64 612 124
rect 554 50 612 64
rect 642 150 700 158
rect 642 72 654 150
rect 688 72 700 150
rect 642 50 700 72
rect 730 120 788 158
rect 730 60 742 120
rect 776 60 788 120
rect 730 50 788 60
rect 818 150 876 158
rect 818 72 830 150
rect 864 72 876 150
rect 818 50 876 72
rect 906 120 964 158
rect 906 60 918 120
rect 952 60 964 120
rect 906 50 964 60
rect 994 150 1052 158
rect 994 72 1006 150
rect 1040 72 1052 150
rect 994 50 1052 72
rect 1082 118 1140 158
rect 1082 58 1094 118
rect 1128 58 1140 118
rect 1082 50 1140 58
rect 1170 150 1230 158
rect 1170 72 1182 150
rect 1216 72 1230 150
rect 1170 50 1230 72
rect 1260 118 1318 158
rect 1260 58 1272 118
rect 1306 58 1318 118
rect 1260 50 1318 58
rect 1348 150 1406 158
rect 1348 72 1360 150
rect 1394 72 1406 150
rect 1348 50 1406 72
<< pdiff >>
rect 28 480 81 496
rect 28 394 36 480
rect 70 394 81 480
rect 28 352 81 394
rect 111 476 168 496
rect 111 360 122 476
rect 156 360 168 476
rect 111 352 168 360
rect 198 482 256 496
rect 198 407 210 482
rect 244 407 256 482
rect 198 352 256 407
rect 286 476 344 496
rect 286 360 298 476
rect 332 360 344 476
rect 286 352 344 360
rect 374 484 432 496
rect 374 408 386 484
rect 420 408 432 484
rect 374 352 432 408
rect 462 476 524 496
rect 462 368 478 476
rect 512 368 524 476
rect 462 352 524 368
rect 554 484 612 496
rect 554 409 566 484
rect 600 409 612 484
rect 554 352 612 409
rect 642 476 700 496
rect 642 368 654 476
rect 688 368 700 476
rect 642 352 700 368
rect 730 484 788 496
rect 730 409 742 484
rect 776 409 788 484
rect 730 352 788 409
rect 818 476 876 496
rect 818 368 830 476
rect 864 368 876 476
rect 818 352 876 368
rect 906 484 964 496
rect 906 409 918 484
rect 952 409 964 484
rect 906 352 964 409
rect 994 476 1052 496
rect 994 368 1006 476
rect 1040 368 1052 476
rect 994 352 1052 368
rect 1082 484 1140 496
rect 1082 409 1094 484
rect 1128 409 1140 484
rect 1082 352 1140 409
rect 1170 476 1230 496
rect 1170 368 1184 476
rect 1218 368 1230 476
rect 1170 352 1230 368
rect 1260 484 1318 496
rect 1260 409 1272 484
rect 1306 409 1318 484
rect 1260 352 1318 409
rect 1348 476 1406 496
rect 1348 368 1360 476
rect 1394 368 1406 476
rect 1348 352 1406 368
<< ndiffc >>
rect 36 64 70 132
rect 122 72 156 150
rect 210 64 244 124
rect 298 72 332 150
rect 386 64 420 124
rect 478 72 512 150
rect 566 64 600 124
rect 654 72 688 150
rect 742 60 776 120
rect 830 72 864 150
rect 918 60 952 120
rect 1006 72 1040 150
rect 1094 58 1128 118
rect 1182 72 1216 150
rect 1272 58 1306 118
rect 1360 72 1394 150
<< pdiffc >>
rect 36 394 70 480
rect 122 360 156 476
rect 210 407 244 482
rect 298 360 332 476
rect 386 408 420 484
rect 478 368 512 476
rect 566 409 600 484
rect 654 368 688 476
rect 742 409 776 484
rect 830 368 864 476
rect 918 409 952 484
rect 1006 368 1040 476
rect 1094 409 1128 484
rect 1184 368 1218 476
rect 1272 409 1306 484
rect 1360 368 1394 476
<< poly >>
rect 81 496 111 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 524 496 554 522
rect 612 496 642 522
rect 700 496 730 522
rect 788 496 818 522
rect 876 496 906 522
rect 964 496 994 522
rect 1052 496 1082 522
rect 1140 496 1170 522
rect 1230 496 1260 522
rect 1318 496 1348 522
rect 81 288 111 352
rect 168 288 198 352
rect 256 288 286 352
rect 344 288 374 352
rect 44 278 374 288
rect 432 290 462 352
rect 524 290 554 352
rect 612 290 642 352
rect 700 290 730 352
rect 788 290 818 352
rect 876 290 906 352
rect 964 290 994 352
rect 1052 290 1082 352
rect 1140 290 1170 352
rect 1230 290 1260 352
rect 1318 290 1348 352
rect 432 280 1366 290
rect 44 244 60 278
rect 360 244 376 278
rect 432 246 456 280
rect 1328 246 1382 280
rect 44 234 374 244
rect 81 158 111 234
rect 168 158 198 234
rect 256 158 286 234
rect 344 158 374 234
rect 432 234 1366 246
rect 432 158 462 234
rect 524 158 554 234
rect 612 158 642 234
rect 700 158 730 234
rect 788 158 818 234
rect 876 158 906 234
rect 964 158 994 234
rect 1052 158 1082 234
rect 1140 158 1170 234
rect 1230 158 1260 234
rect 1318 158 1348 234
rect 81 24 111 50
rect 168 24 198 50
rect 256 24 286 50
rect 344 24 374 50
rect 432 24 462 50
rect 524 24 554 50
rect 612 24 642 50
rect 700 24 730 50
rect 788 24 818 50
rect 876 24 906 50
rect 964 24 994 50
rect 1052 24 1082 50
rect 1140 24 1170 50
rect 1230 24 1260 50
rect 1318 24 1348 50
<< polycont >>
rect 60 244 360 278
rect 456 246 1328 280
<< locali >>
rect 0 561 1472 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 526 1472 527
rect 36 480 70 526
rect 36 378 70 394
rect 122 476 156 492
rect 210 482 244 526
rect 210 391 244 407
rect 298 476 332 492
rect 122 357 156 360
rect 386 484 420 526
rect 386 392 420 408
rect 478 476 512 492
rect 298 357 332 360
rect 566 484 600 526
rect 566 393 600 409
rect 654 476 688 492
rect 478 359 512 368
rect 742 484 776 526
rect 742 393 776 409
rect 830 476 864 492
rect 654 359 688 368
rect 918 484 952 526
rect 918 393 952 409
rect 1006 476 1040 492
rect 830 359 864 368
rect 1094 484 1128 526
rect 1094 393 1128 409
rect 1184 476 1218 492
rect 1006 359 1040 368
rect 1272 484 1306 526
rect 1272 393 1306 409
rect 1360 476 1394 492
rect 1184 359 1218 368
rect 1360 359 1394 368
rect 122 323 444 357
rect 478 325 1444 359
rect 410 291 444 323
rect 38 278 376 289
rect 38 244 60 278
rect 360 244 376 278
rect 410 280 1344 291
rect 410 246 456 280
rect 1328 246 1344 280
rect 410 210 444 246
rect 122 174 444 210
rect 1378 208 1444 325
rect 478 174 1444 208
rect 122 150 156 174
rect 36 132 70 148
rect 36 21 70 64
rect 298 150 332 174
rect 122 56 156 72
rect 210 124 244 140
rect 210 21 244 64
rect 478 150 512 174
rect 298 56 332 72
rect 386 124 420 140
rect 386 21 420 64
rect 654 150 688 174
rect 478 56 512 72
rect 566 124 600 140
rect 566 21 600 64
rect 830 150 864 174
rect 654 56 688 72
rect 742 120 776 140
rect 742 21 776 60
rect 1006 150 1040 174
rect 830 56 864 72
rect 918 120 952 140
rect 918 21 952 60
rect 1182 150 1216 174
rect 1006 56 1040 72
rect 1094 118 1128 140
rect 1094 21 1128 58
rect 1360 150 1394 174
rect 1182 56 1216 72
rect 1272 118 1306 140
rect 1272 21 1306 58
rect 1360 56 1394 72
rect 0 17 1472 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_11
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 170 255 204 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 187 272 187 272 0 FreeSans 200 0 0 0 A
flabel locali s 255 255 289 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 272 272 272 272 0 FreeSans 200 0 0 0 A
flabel locali s 68 255 102 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 1394 306 1428 340 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 1411 323 1411 323 0 FreeSans 200 0 0 0 Y
flabel locali s 1394 187 1428 221 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 1411 204 1411 204 0 FreeSans 200 0 0 0 Y
flabel locali s 85 272 85 272 0 FreeSans 200 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_11.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
