magic
tech sky130A
magscale 1 2
timestamp 1740499863
<< nwell >>
rect -38 262 2430 582
<< pwell >>
rect 0 34 2392 204
rect 0 32 1656 34
rect 2022 32 2300 34
rect 0 24 1472 32
rect 0 22 736 24
rect 1099 22 1104 24
rect 26 -20 90 22
<< pmos >>
rect 112 298 142 496
rect 224 412 276 496
rect 442 298 472 496
rect 528 298 558 496
rect 752 298 782 496
rect 856 298 886 496
rect 948 298 978 496
rect 1200 298 1230 496
rect 1396 298 1426 496
rect 1592 298 1622 496
rect 1698 298 1728 496
rect 1784 298 1814 496
rect 2012 298 2042 496
rect 2098 298 2128 496
rect 2212 298 2242 496
<< nmoslvt >>
rect 112 48 142 178
rect 224 48 276 178
rect 442 48 472 178
rect 528 48 558 178
rect 752 48 782 178
rect 856 48 886 178
rect 948 48 978 178
rect 1200 48 1230 178
rect 1300 48 1330 178
rect 1520 48 1550 178
rect 1698 48 1728 178
rect 1784 48 1814 178
rect 2012 48 2042 178
rect 2098 48 2128 178
rect 2212 48 2242 178
<< ndiff >>
rect 27 166 112 178
rect 27 132 35 166
rect 69 132 112 166
rect 27 48 112 132
rect 142 90 224 178
rect 142 56 168 90
rect 202 56 224 90
rect 142 48 224 56
rect 276 166 330 178
rect 276 132 288 166
rect 322 132 330 166
rect 276 48 330 132
rect 384 166 442 178
rect 384 132 397 166
rect 431 132 442 166
rect 384 48 442 132
rect 472 90 528 178
rect 472 56 483 90
rect 517 56 528 90
rect 472 48 528 56
rect 558 166 634 178
rect 558 132 592 166
rect 626 132 634 166
rect 558 48 634 132
rect 698 94 752 178
rect 698 60 707 94
rect 741 60 752 94
rect 698 48 752 60
rect 782 170 856 178
rect 782 136 793 170
rect 827 136 856 170
rect 782 48 856 136
rect 886 94 948 178
rect 886 60 897 94
rect 931 60 948 94
rect 886 48 948 60
rect 978 166 1068 178
rect 978 132 1026 166
rect 1060 132 1068 166
rect 978 48 1068 132
rect 1146 94 1200 178
rect 1146 60 1155 94
rect 1189 60 1200 94
rect 1146 48 1200 60
rect 1230 166 1300 178
rect 1230 132 1241 166
rect 1275 132 1300 166
rect 1230 48 1300 132
rect 1330 164 1520 178
rect 1330 130 1474 164
rect 1508 130 1520 164
rect 1330 48 1520 130
rect 1550 48 1698 178
rect 1728 94 1784 178
rect 1728 60 1739 94
rect 1773 60 1784 94
rect 1728 48 1784 60
rect 1814 164 1904 178
rect 1814 130 1862 164
rect 1896 130 1904 164
rect 1814 48 1904 130
rect 1958 164 2012 178
rect 1958 130 1967 164
rect 2001 130 2012 164
rect 1958 48 2012 130
rect 2042 92 2098 178
rect 2042 58 2053 92
rect 2087 58 2098 92
rect 2042 48 2098 58
rect 2128 164 2212 178
rect 2128 130 2164 164
rect 2198 130 2212 164
rect 2128 48 2212 130
rect 2242 170 2322 178
rect 2242 56 2256 170
rect 2290 56 2322 170
rect 2242 48 2322 56
<< pdiff >>
rect 27 476 112 496
rect 27 310 35 476
rect 69 310 112 476
rect 27 298 112 310
rect 142 488 224 496
rect 142 420 162 488
rect 196 420 224 488
rect 142 412 224 420
rect 276 476 330 496
rect 276 424 288 476
rect 322 424 330 476
rect 276 412 330 424
rect 384 476 442 496
rect 142 298 192 412
rect 384 306 397 476
rect 431 306 442 476
rect 384 298 442 306
rect 472 482 528 496
rect 472 424 483 482
rect 517 424 528 482
rect 472 298 528 424
rect 558 476 634 496
rect 558 310 592 476
rect 626 310 634 476
rect 558 298 634 310
rect 698 476 752 496
rect 698 322 707 476
rect 741 322 752 476
rect 698 298 752 322
rect 782 298 856 496
rect 886 480 948 496
rect 886 426 897 480
rect 931 426 948 480
rect 886 298 948 426
rect 978 470 1068 496
rect 978 312 1026 470
rect 1060 312 1068 470
rect 978 298 1068 312
rect 1146 484 1200 496
rect 1146 318 1155 484
rect 1189 318 1200 484
rect 1146 298 1200 318
rect 1230 476 1396 496
rect 1230 306 1241 476
rect 1275 306 1396 476
rect 1230 298 1396 306
rect 1426 476 1592 496
rect 1426 306 1474 476
rect 1508 306 1592 476
rect 1426 298 1592 306
rect 1622 298 1698 496
rect 1728 486 1784 496
rect 1728 452 1739 486
rect 1773 452 1784 486
rect 1728 298 1784 452
rect 1814 476 1904 496
rect 1814 310 1862 476
rect 1896 310 1904 476
rect 1814 298 1904 310
rect 1958 476 2012 496
rect 1958 310 1967 476
rect 2001 310 2012 476
rect 1958 298 2012 310
rect 2042 478 2098 496
rect 2042 318 2053 478
rect 2087 318 2098 478
rect 2042 298 2098 318
rect 2128 476 2212 496
rect 2128 310 2164 476
rect 2198 310 2212 476
rect 2128 298 2212 310
rect 2242 488 2322 496
rect 2242 306 2256 488
rect 2290 306 2322 488
rect 2242 298 2322 306
<< ndiffc >>
rect 35 132 69 166
rect 168 56 202 90
rect 288 132 322 166
rect 397 132 431 166
rect 483 56 517 90
rect 592 132 626 166
rect 707 60 741 94
rect 793 136 827 170
rect 897 60 931 94
rect 1026 132 1060 166
rect 1155 60 1189 94
rect 1241 132 1275 166
rect 1474 130 1508 164
rect 1739 60 1773 94
rect 1862 130 1896 164
rect 1967 130 2001 164
rect 2053 58 2087 92
rect 2164 130 2198 164
rect 2256 56 2290 170
<< pdiffc >>
rect 35 310 69 476
rect 162 420 196 488
rect 288 424 322 476
rect 397 306 431 476
rect 483 424 517 482
rect 592 310 626 476
rect 707 322 741 476
rect 897 426 931 480
rect 1026 312 1060 470
rect 1155 318 1189 484
rect 1241 306 1275 476
rect 1474 306 1508 476
rect 1739 452 1773 486
rect 1862 310 1896 476
rect 1967 310 2001 476
rect 2053 318 2087 478
rect 2164 310 2198 476
rect 2256 306 2290 488
<< poly >>
rect 112 496 142 522
rect 224 496 276 522
rect 442 496 472 522
rect 528 496 558 522
rect 752 496 782 522
rect 856 496 886 522
rect 948 496 978 522
rect 1200 496 1230 522
rect 1396 496 1426 522
rect 1592 496 1622 522
rect 1698 496 1728 522
rect 1784 496 1814 522
rect 2012 496 2042 522
rect 2098 496 2128 522
rect 2212 496 2242 522
rect 112 266 142 298
rect 224 266 276 412
rect 104 250 158 266
rect 104 216 114 250
rect 148 216 158 250
rect 104 196 158 216
rect 200 250 276 266
rect 200 216 210 250
rect 244 216 276 250
rect 200 196 276 216
rect 318 250 372 266
rect 442 250 472 298
rect 528 268 558 298
rect 318 216 328 250
rect 362 216 472 250
rect 318 196 372 216
rect 112 178 142 196
rect 224 178 276 196
rect 442 178 472 216
rect 514 250 568 268
rect 514 216 524 250
rect 558 216 568 250
rect 514 198 568 216
rect 624 250 678 268
rect 752 250 782 298
rect 856 266 886 298
rect 948 266 978 298
rect 1200 266 1230 298
rect 1396 266 1426 298
rect 1592 266 1622 298
rect 1698 266 1728 298
rect 1784 266 1814 298
rect 624 216 634 250
rect 668 216 782 250
rect 624 198 678 216
rect 528 178 558 198
rect 752 178 782 216
rect 852 250 906 266
rect 852 216 862 250
rect 896 216 906 250
rect 852 196 906 216
rect 948 250 1002 266
rect 948 216 958 250
rect 992 216 1002 250
rect 948 196 1002 216
rect 1132 250 1230 266
rect 1132 216 1142 250
rect 1176 216 1230 250
rect 1132 196 1230 216
rect 856 178 886 196
rect 948 178 978 196
rect 1200 178 1230 196
rect 1300 250 1354 266
rect 1300 216 1310 250
rect 1344 216 1354 250
rect 1300 196 1354 216
rect 1396 250 1450 266
rect 1396 216 1406 250
rect 1440 226 1450 250
rect 1592 250 1646 266
rect 1440 216 1550 226
rect 1396 196 1550 216
rect 1592 216 1602 250
rect 1636 216 1646 250
rect 1592 196 1646 216
rect 1688 250 1742 266
rect 1688 216 1698 250
rect 1732 216 1742 250
rect 1688 196 1742 216
rect 1784 250 1838 266
rect 1784 216 1794 250
rect 1828 216 1838 250
rect 1784 196 1838 216
rect 1880 250 1938 268
rect 1880 216 1890 250
rect 1924 246 1938 250
rect 2012 246 2042 298
rect 2098 268 2128 298
rect 1924 216 2042 246
rect 1880 212 2042 216
rect 1880 198 1938 212
rect 1300 178 1330 196
rect 1520 178 1550 196
rect 1698 178 1728 196
rect 1784 178 1814 196
rect 2012 178 2042 212
rect 2084 250 2142 268
rect 2212 250 2242 298
rect 2084 216 2096 250
rect 2130 216 2242 250
rect 2084 198 2142 216
rect 2098 178 2128 198
rect 2212 178 2242 216
rect 112 22 142 48
rect 224 22 276 48
rect 442 22 472 48
rect 528 22 558 48
rect 752 22 782 48
rect 856 22 886 48
rect 948 22 978 48
rect 1200 22 1230 48
rect 1300 22 1330 48
rect 1520 22 1550 48
rect 1698 22 1728 48
rect 1784 22 1814 48
rect 2012 22 2042 48
rect 2098 22 2128 48
rect 2212 22 2242 48
<< polycont >>
rect 114 216 148 250
rect 210 216 244 250
rect 328 216 362 250
rect 524 216 558 250
rect 634 216 668 250
rect 862 216 896 250
rect 958 216 992 250
rect 1142 216 1176 250
rect 1310 216 1344 250
rect 1406 216 1440 250
rect 1602 216 1636 250
rect 1698 216 1732 250
rect 1794 216 1828 250
rect 1890 216 1924 250
rect 2096 216 2130 250
<< locali >>
rect 0 561 2392 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 526 2392 527
rect 35 476 69 492
rect 162 488 196 526
rect 162 314 196 420
rect 288 476 322 492
rect 35 166 69 310
rect 288 266 322 424
rect 397 476 431 492
rect 483 482 517 526
rect 483 408 517 424
rect 592 476 626 492
rect 104 250 158 266
rect 104 216 114 250
rect 148 216 158 250
rect 104 196 158 216
rect 210 250 244 266
rect 210 162 244 216
rect 69 132 210 162
rect 35 128 210 132
rect 288 250 362 266
rect 288 216 328 250
rect 288 196 362 216
rect 397 250 431 306
rect 592 268 626 310
rect 707 476 741 492
rect 897 480 931 526
rect 897 408 931 426
rect 1026 470 1060 492
rect 741 322 992 340
rect 707 306 992 322
rect 524 250 558 268
rect 397 216 524 250
rect 288 166 322 196
rect 35 116 69 128
rect 288 116 322 132
rect 397 166 431 216
rect 524 198 558 216
rect 592 250 678 268
rect 592 216 634 250
rect 668 216 678 250
rect 592 198 678 216
rect 397 116 431 132
rect 592 166 626 198
rect 592 116 626 132
rect 793 170 827 306
rect 862 250 896 266
rect 862 196 896 216
rect 958 250 992 306
rect 958 196 992 216
rect 793 120 827 136
rect 1026 166 1060 312
rect 1155 484 1189 526
rect 1155 302 1189 318
rect 1241 476 1275 492
rect 1132 250 1186 266
rect 1132 216 1142 250
rect 1176 216 1186 250
rect 1132 196 1186 216
rect 1026 116 1060 132
rect 1241 166 1275 306
rect 1474 476 1508 492
rect 1739 486 1773 526
rect 1739 436 1773 452
rect 1862 476 1896 492
rect 1310 250 1344 266
rect 1310 196 1344 216
rect 1406 250 1440 266
rect 1406 196 1440 216
rect 1241 114 1275 132
rect 1474 164 1508 306
rect 1698 320 1862 354
rect 1602 250 1636 266
rect 1602 196 1636 216
rect 1698 250 1732 320
rect 1862 268 1896 310
rect 1967 476 2001 492
rect 1698 196 1732 216
rect 1794 250 1828 266
rect 1794 162 1828 216
rect 1508 130 1828 162
rect 1474 128 1828 130
rect 1862 250 1924 268
rect 1862 216 1890 250
rect 1862 198 1924 216
rect 1967 250 2001 310
rect 2053 478 2087 526
rect 2053 302 2087 318
rect 2164 476 2198 492
rect 2164 308 2198 310
rect 2256 488 2290 526
rect 2084 250 2130 268
rect 1967 216 2096 250
rect 1862 164 1896 198
rect 1474 114 1508 128
rect 1862 114 1896 130
rect 1967 164 2001 216
rect 2084 198 2130 216
rect 1967 114 2001 130
rect 2164 164 2218 308
rect 2256 290 2290 306
rect 2256 170 2290 186
rect 2164 114 2198 130
rect 152 56 168 90
rect 202 56 218 90
rect 466 56 483 90
rect 517 56 534 90
rect 690 60 707 94
rect 741 60 758 94
rect 880 60 897 94
rect 931 60 948 94
rect 1138 60 1155 94
rect 1189 60 1206 94
rect 1722 60 1739 94
rect 1773 60 1790 94
rect 2053 92 2087 108
rect 168 21 202 56
rect 483 21 517 56
rect 707 21 741 60
rect 897 21 931 60
rect 1155 21 1189 60
rect 1739 21 1773 60
rect 2053 21 2087 58
rect 2256 21 2290 56
rect 0 17 2392 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 210 128 244 162
rect 862 216 896 250
rect 1026 132 1060 166
rect 1310 216 1344 250
rect 1406 216 1440 250
rect 1602 216 1636 250
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 1290 442 1636 444
rect 862 408 1636 442
rect 862 262 896 408
rect 856 250 902 262
rect 1310 258 1344 408
rect 1602 266 1636 408
rect 856 216 862 250
rect 896 216 902 250
rect 856 196 902 216
rect 1304 250 1350 258
rect 1304 216 1310 250
rect 1344 216 1350 250
rect 1304 204 1350 216
rect 1400 250 1446 264
rect 1400 216 1406 250
rect 1440 216 1446 250
rect 1400 210 1446 216
rect 1594 250 1644 266
rect 1594 216 1602 250
rect 1636 216 1644 250
rect 198 162 276 168
rect 862 162 896 196
rect 198 128 210 162
rect 244 128 896 162
rect 1020 166 1066 178
rect 1020 132 1026 166
rect 1060 132 1066 166
rect 198 122 276 128
rect 1020 120 1066 132
rect 1406 120 1440 210
rect 1594 204 1644 216
rect 1020 86 1440 120
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
rlabel comment s 0 0 0 0 4 pulsed_dfxtp_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 2392 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 119 221 153 255 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel locali s 136 238 136 238 0 FreeSans 200 0 0 0 CLK
flabel locali 1150 221 1184 255 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali 1167 238 1167 238 0 FreeSans 200 0 0 0 D
flabel locali 2170 221 2204 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali 2185 228 2185 238 0 FreeSans 200 0 0 0 Q
<< properties >>
string FIXED_BBOX 0 0 2392 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
