magic
tech sky130A
magscale 1 2
timestamp 1739976054
<< nwell >>
rect -38 262 1142 582
<< pwell >>
rect 0 30 1104 204
rect 0 28 920 30
rect 26 -22 68 28
rect 276 22 736 28
rect 302 -20 366 22
<< pmos >>
rect 166 298 196 496
rect 356 298 386 496
rect 442 298 472 496
rect 528 298 558 496
rect 718 298 748 496
rect 804 298 834 496
rect 890 298 920 496
rect 976 298 1006 496
<< nmoslvt >>
rect 166 48 196 178
rect 356 48 386 178
rect 442 48 472 178
rect 528 48 558 178
rect 718 48 748 178
rect 804 48 834 178
rect 890 48 920 178
rect 976 48 1006 178
<< ndiff >>
rect 27 150 166 178
rect 27 56 40 150
rect 155 56 166 150
rect 27 48 166 56
rect 196 166 249 178
rect 196 72 207 166
rect 241 72 249 166
rect 196 48 249 72
rect 303 105 356 178
rect 303 71 311 105
rect 345 71 356 105
rect 303 48 356 71
rect 386 48 442 178
rect 472 90 528 178
rect 472 56 483 90
rect 517 56 528 90
rect 472 48 528 56
rect 558 150 611 178
rect 558 72 569 150
rect 603 72 611 150
rect 558 48 611 72
rect 665 94 718 178
rect 665 60 673 94
rect 707 60 718 94
rect 665 48 718 60
rect 748 170 804 178
rect 748 72 759 170
rect 793 72 804 170
rect 748 48 804 72
rect 834 132 890 178
rect 834 56 845 132
rect 879 56 890 132
rect 834 48 890 56
rect 920 170 976 178
rect 920 72 931 170
rect 965 72 976 170
rect 920 48 976 72
rect 1006 170 1077 178
rect 1006 56 1017 170
rect 1051 56 1077 170
rect 1006 48 1077 56
<< pdiff >>
rect 27 476 166 496
rect 27 316 36 476
rect 155 316 166 476
rect 27 298 166 316
rect 196 476 249 496
rect 196 310 207 476
rect 241 310 249 476
rect 196 298 249 310
rect 303 476 356 496
rect 303 316 311 476
rect 345 316 356 476
rect 303 298 356 316
rect 386 488 442 496
rect 386 454 397 488
rect 431 454 442 488
rect 386 298 442 454
rect 472 476 528 496
rect 472 316 483 476
rect 517 316 528 476
rect 472 298 528 316
rect 558 476 611 496
rect 558 332 569 476
rect 603 332 611 476
rect 558 298 611 332
rect 665 484 718 496
rect 665 388 673 484
rect 707 388 718 484
rect 665 298 718 388
rect 748 476 804 496
rect 748 306 759 476
rect 793 306 804 476
rect 748 298 804 306
rect 834 488 890 496
rect 834 338 845 488
rect 879 338 890 488
rect 834 298 890 338
rect 920 476 976 496
rect 920 306 931 476
rect 965 306 976 476
rect 920 298 976 306
rect 1006 488 1077 496
rect 1006 306 1017 488
rect 1051 306 1077 488
rect 1006 298 1077 306
<< ndiffc >>
rect 40 56 155 150
rect 207 72 241 166
rect 311 71 345 105
rect 483 56 517 90
rect 569 72 603 150
rect 673 60 707 94
rect 759 72 793 170
rect 845 56 879 132
rect 931 72 965 170
rect 1017 56 1051 170
<< pdiffc >>
rect 36 316 155 476
rect 207 310 241 476
rect 311 316 345 476
rect 397 454 431 488
rect 483 316 517 476
rect 569 332 603 476
rect 673 388 707 484
rect 759 306 793 476
rect 845 338 879 488
rect 931 306 965 476
rect 1017 306 1051 488
<< poly >>
rect 166 496 196 522
rect 356 496 386 522
rect 442 496 472 522
rect 528 496 558 522
rect 718 496 748 522
rect 804 496 834 522
rect 890 496 920 522
rect 976 496 1006 522
rect 166 266 196 298
rect 356 266 386 298
rect 442 266 472 298
rect 528 266 558 298
rect 718 266 748 298
rect 804 266 834 298
rect 122 250 196 266
rect 122 216 134 250
rect 168 216 196 250
rect 122 200 196 216
rect 316 250 386 266
rect 316 216 328 250
rect 362 216 386 250
rect 316 200 386 216
rect 428 250 482 266
rect 428 216 438 250
rect 472 216 482 250
rect 428 200 482 216
rect 524 250 578 266
rect 524 216 534 250
rect 568 216 578 250
rect 524 200 578 216
rect 670 250 834 266
rect 670 216 686 250
rect 720 246 834 250
rect 890 262 920 298
rect 976 262 1006 298
rect 890 246 1006 262
rect 720 230 1006 246
rect 720 216 920 230
rect 670 200 920 216
rect 166 178 196 200
rect 356 178 386 200
rect 442 178 472 200
rect 528 178 558 200
rect 718 178 748 200
rect 804 178 834 200
rect 890 178 920 200
rect 976 178 1006 230
rect 166 22 196 48
rect 356 22 386 48
rect 442 22 472 48
rect 528 22 558 48
rect 718 22 748 48
rect 804 22 834 48
rect 890 22 920 48
rect 976 22 1006 48
<< polycont >>
rect 134 216 168 250
rect 328 216 362 250
rect 438 216 472 250
rect 534 216 568 250
rect 686 216 720 250
<< locali >>
rect 0 561 1104 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 526 1104 527
rect 34 476 155 526
rect 34 316 36 476
rect 34 300 155 316
rect 207 476 241 492
rect 82 250 172 266
rect 82 216 134 250
rect 168 216 172 250
rect 82 200 172 216
rect 207 240 241 310
rect 311 476 345 492
rect 397 488 431 526
rect 397 438 431 454
rect 483 476 517 492
rect 345 370 483 404
rect 311 300 345 316
rect 398 266 448 336
rect 569 476 603 492
rect 673 484 707 526
rect 673 372 707 388
rect 759 476 793 492
rect 603 332 646 350
rect 569 316 646 332
rect 483 300 517 316
rect 612 266 646 316
rect 845 488 879 526
rect 845 322 879 338
rect 931 476 965 492
rect 759 298 793 306
rect 314 250 364 266
rect 314 240 328 250
rect 207 216 328 240
rect 362 216 364 250
rect 207 200 364 216
rect 398 250 476 266
rect 398 216 438 250
rect 472 216 476 250
rect 398 200 476 216
rect 524 250 578 266
rect 524 216 534 250
rect 568 216 578 250
rect 524 200 578 216
rect 612 250 724 266
rect 612 216 686 250
rect 720 216 724 250
rect 612 200 724 216
rect 759 260 820 298
rect 931 260 965 306
rect 1017 488 1051 526
rect 1017 288 1051 306
rect 759 208 965 260
rect 207 166 241 200
rect 612 166 646 200
rect 36 150 155 166
rect 36 56 40 150
rect 398 150 646 166
rect 398 132 569 150
rect 207 56 241 72
rect 311 105 345 121
rect 398 89 432 132
rect 345 71 432 89
rect 36 21 155 56
rect 311 55 432 71
rect 466 90 534 98
rect 466 56 483 90
rect 517 56 534 90
rect 603 132 646 150
rect 759 172 820 208
rect 759 170 793 172
rect 569 56 603 72
rect 673 94 707 110
rect 483 21 518 56
rect 673 21 707 60
rect 931 170 965 208
rect 759 56 793 72
rect 845 132 879 148
rect 931 56 965 72
rect 1017 170 1051 186
rect 845 21 879 56
rect 1017 21 1051 56
rect 0 17 1104 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ao21b_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 136 221 170 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 153 238 153 238 0 FreeSans 200 0 0 0 A
flabel locali s 429 221 463 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 446 238 446 238 0 FreeSans 200 0 0 0 B
flabel locali s 531 221 565 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 548 238 548 238 0 FreeSans 200 0 0 0 C
flabel locali s 769 221 803 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 786 238 786 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__ao21b_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1104 220
string MASKHINTS_NSDM 0 -38 1104 209
string MASKHINTS_PSDM 0 273 1104 582
<< end >>
