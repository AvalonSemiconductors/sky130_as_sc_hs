VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.605 2.050 0.775 2.630 ;
        RECT 1.490 1.910 1.660 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.700 ;
        RECT 1.490 0.105 1.660 0.760 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.210 1.810 1.020 ;
        RECT 0.110 -0.100 0.450 0.210 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.210 0.450 1.540 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.910 1.320 2.420 ;
        RECT 1.150 1.460 1.320 1.910 ;
        RECT 1.150 1.260 1.385 1.460 ;
        RECT 1.150 0.800 1.320 1.260 ;
        RECT 1.050 0.290 1.320 0.800 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.170 1.880 0.340 2.420 ;
        RECT 0.170 1.710 0.880 1.880 ;
        RECT 0.710 1.560 0.880 1.710 ;
        RECT 0.710 1.230 0.980 1.560 ;
        RECT 0.710 1.040 0.880 1.230 ;
        RECT 0.175 0.870 0.880 1.040 ;
        RECT 0.175 0.290 0.345 0.870 ;
  END
END sky130_as_sc_hs__buff_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_11
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.180 1.890 0.350 2.630 ;
        RECT 1.050 1.955 1.220 2.630 ;
        RECT 1.930 1.960 2.100 2.630 ;
        RECT 2.830 1.965 3.000 2.630 ;
        RECT 3.710 1.965 3.880 2.630 ;
        RECT 4.590 1.965 4.760 2.630 ;
        RECT 5.470 1.965 5.640 2.630 ;
        RECT 6.360 1.965 6.530 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.105 0.350 0.740 ;
        RECT 1.050 0.105 1.220 0.700 ;
        RECT 1.930 0.105 2.100 0.700 ;
        RECT 2.830 0.105 3.000 0.700 ;
        RECT 3.710 0.105 3.880 0.700 ;
        RECT 4.590 0.105 4.760 0.700 ;
        RECT 5.470 0.105 5.640 0.700 ;
        RECT 6.360 0.105 6.530 0.700 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 7.120 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 1.220 1.880 1.445 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.230200 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.795 2.560 2.460 ;
        RECT 3.270 1.795 3.440 2.460 ;
        RECT 4.150 1.795 4.320 2.460 ;
        RECT 5.030 1.795 5.200 2.460 ;
        RECT 5.920 1.795 6.090 2.460 ;
        RECT 6.800 1.795 6.970 2.460 ;
        RECT 7.140 1.795 7.330 1.870 ;
        RECT 2.390 1.625 7.330 1.795 ;
        RECT 7.080 1.040 7.330 1.625 ;
        RECT 2.390 0.870 7.330 1.040 ;
        RECT 2.390 0.280 2.560 0.870 ;
        RECT 3.270 0.280 3.440 0.870 ;
        RECT 4.150 0.280 4.320 0.870 ;
        RECT 5.030 0.280 5.200 0.870 ;
        RECT 5.910 0.280 6.080 0.870 ;
        RECT 6.800 0.280 6.970 0.870 ;
        RECT 7.140 0.700 7.330 0.870 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.610 1.785 0.780 2.460 ;
        RECT 1.490 1.785 1.660 2.460 ;
        RECT 0.610 1.615 2.220 1.785 ;
        RECT 2.050 1.455 2.220 1.615 ;
        RECT 2.050 1.230 6.910 1.455 ;
        RECT 2.050 1.050 2.220 1.230 ;
        RECT 0.610 0.870 2.220 1.050 ;
        RECT 0.610 0.280 0.780 0.870 ;
        RECT 1.490 0.280 1.660 0.870 ;
  END
END sky130_as_sc_hs__buff_11

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_3
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.110 -0.075 0.380 0.220 ;
        RECT 0.110 -0.110 0.360 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.980 0.580 1.580 ;
        RECT 0.140 0.105 1.210 0.980 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.140 1.830 1.210 2.630 ;
        RECT 0.830 1.150 1.170 1.830 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
END sky130_as_sc_hs__decap_3

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.110 0.240 1.730 1.020 ;
        RECT 0.130 0.220 1.600 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.170 1.850 1.670 2.630 ;
        RECT 1.270 1.180 1.610 1.850 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.900 0.580 1.580 ;
        RECT 0.180 0.105 1.660 0.900 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_4

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.220 7.120 1.020 ;
        RECT 0.120 -0.110 0.520 0.220 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.360 1.690 6.980 2.630 ;
        RECT 0.600 1.340 0.850 1.690 ;
        RECT 0.560 1.140 0.890 1.340 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 6.390 0.940 6.720 1.520 ;
        RECT 0.360 0.105 6.970 0.940 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_16

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.850 8.040 1.020 ;
        RECT 0.090 0.260 8.145 0.850 ;
        RECT 0.090 0.240 8.040 0.260 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.280 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.620 0.105 0.790 0.640 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.840 ;
        RECT 0.000 -0.085 8.280 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.186000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 1.220 0.440 1.580 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.331250 ;
    PORT
      LAYER li1 ;
        RECT 7.915 1.690 8.085 2.420 ;
        RECT 7.690 1.150 8.085 1.690 ;
        RECT 7.915 0.300 8.085 1.150 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.163500 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.910 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.450 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.180 1.070 1.450 ;
        RECT 0.610 0.980 0.780 1.180 ;
        RECT 1.240 1.010 1.410 1.590 ;
        RECT 0.190 0.810 0.780 0.980 ;
        RECT 1.060 0.840 1.410 1.010 ;
        RECT 0.190 0.280 0.360 0.810 ;
        RECT 1.060 0.280 1.230 0.840 ;
        RECT 2.080 0.280 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 2.420 1.560 2.630 1.890 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.850 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.420 1.050 2.630 1.380 ;
        RECT 2.800 0.880 2.970 1.610 ;
        RECT 4.170 1.520 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.560 5.100 1.890 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 6.670 1.790 6.860 1.850 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 2.710 0.710 2.970 0.880 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 2.710 0.600 2.880 0.710 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 1.050 5.110 1.380 ;
        RECT 5.280 0.880 5.450 1.620 ;
        RECT 6.670 1.520 6.860 1.620 ;
        RECT 7.030 1.590 7.200 2.030 ;
        RECT 6.280 1.230 6.490 1.310 ;
        RECT 7.030 1.260 7.470 1.590 ;
        RECT 7.030 1.230 7.200 1.260 ;
        RECT 5.190 0.710 5.450 0.880 ;
        RECT 5.790 0.830 6.000 1.160 ;
        RECT 6.280 1.060 7.200 1.230 ;
        RECT 6.280 0.980 6.490 1.060 ;
        RECT 7.030 0.790 7.200 1.060 ;
        RECT 5.190 0.600 5.360 0.710 ;
        RECT 5.030 0.430 5.360 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 1.170 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 1.170 1.590 1.470 1.610 ;
        RECT 0.760 1.180 1.070 1.450 ;
        RECT 0.760 0.630 0.900 1.180 ;
        RECT 2.380 1.100 2.690 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.970 1.330 5.110 1.340 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.690 1.100 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.090 5.170 1.150 ;
        RECT 4.970 1.050 5.110 1.090 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.470 0.630 6.000 0.640 ;
        RECT 0.760 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxtp_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__diode_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.220 0.870 1.020 ;
        RECT 0.210 -0.075 0.390 0.220 ;
    END
  END VNB
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.441000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 0.290 0.740 2.450 ;
    END
  END DIODE
END sky130_as_sc_hs__diode_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_4

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.210 0.360 0.450 2.360 ;
  END
END sky130_as_sc_hs__fill_8

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.730 2.020 0.970 2.260 ;
        RECT 0.490 1.780 1.210 2.020 ;
        RECT 0.490 1.300 0.730 1.780 ;
        RECT 0.970 1.300 1.210 1.780 ;
        RECT 1.690 1.540 1.930 2.260 ;
        RECT 3.130 1.540 3.370 2.260 ;
        RECT 4.090 2.020 4.330 2.260 ;
        RECT 1.690 1.300 2.170 1.540 ;
        RECT 0.490 1.060 1.210 1.300 ;
        RECT 0.250 0.820 0.730 1.060 ;
        RECT 0.970 0.820 1.450 1.060 ;
        RECT 0.250 0.340 0.490 0.820 ;
        RECT 1.210 0.340 1.450 0.820 ;
        RECT 1.930 0.820 2.170 1.300 ;
        RECT 2.410 0.820 2.650 1.540 ;
        RECT 2.890 1.300 3.370 1.540 ;
        RECT 3.850 1.780 4.570 2.020 ;
        RECT 3.850 1.300 4.090 1.780 ;
        RECT 4.330 1.300 4.570 1.780 ;
        RECT 5.050 1.540 5.290 2.260 ;
        RECT 6.490 1.540 6.730 2.260 ;
        RECT 5.050 1.300 5.530 1.540 ;
        RECT 2.890 0.820 3.130 1.300 ;
        RECT 3.850 1.060 4.570 1.300 ;
        RECT 1.930 0.580 3.130 0.820 ;
        RECT 3.610 0.820 4.090 1.060 ;
        RECT 4.330 0.820 4.810 1.060 ;
        RECT 2.170 0.340 2.410 0.580 ;
        RECT 2.650 0.340 2.890 0.580 ;
        RECT 3.610 0.340 3.850 0.820 ;
        RECT 4.570 0.340 4.810 0.820 ;
        RECT 5.290 0.820 5.530 1.300 ;
        RECT 5.770 0.820 6.010 1.540 ;
        RECT 6.250 1.300 6.730 1.540 ;
        RECT 6.250 0.820 6.490 1.300 ;
        RECT 5.290 0.580 6.490 0.820 ;
        RECT 5.530 0.340 5.770 0.580 ;
        RECT 6.010 0.340 6.250 0.580 ;
  END
END sky130_as_sc_hs__fill_16

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.220 1.600 1.020 ;
        RECT 0.120 -0.075 0.380 0.220 ;
        RECT 0.120 -0.110 0.350 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.320 1.610 0.570 2.630 ;
        RECT 1.320 1.610 1.570 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.310 0.105 0.560 0.950 ;
        RECT 1.280 0.280 1.550 0.950 ;
        RECT 1.280 0.105 1.530 0.280 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.624000 ;
    PORT
      LAYER li1 ;
        RECT 0.300 1.120 0.630 1.440 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.468000 ;
    PORT
      LAYER li1 ;
        RECT 0.820 0.310 1.070 2.430 ;
    END
  END Y
END sky130_as_sc_hs__inv_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand2_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.080 1.310 1.020 ;
        RECT 0.210 -0.075 0.380 0.080 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.140 1.610 0.310 2.630 ;
        RECT 1.010 1.640 1.180 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.105 0.310 0.860 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.240750 ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.090 1.190 1.420 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.240750 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.080 0.405 1.420 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.448075 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.040 0.745 2.450 ;
        RECT 0.575 0.920 0.765 1.040 ;
        RECT 0.575 0.750 1.180 0.920 ;
        RECT 1.010 0.360 1.180 0.750 ;
    END
  END Y
END sky130_as_sc_hs__nand2_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.090 1.380 1.020 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.175 1.610 0.345 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.860 ;
        RECT 1.035 0.105 1.205 0.920 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.090 1.205 1.430 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.237000 ;
    PORT
      LAYER li1 ;
        RECT 0.165 1.080 0.435 1.420 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.428675 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.780 1.205 2.460 ;
        RECT 0.605 1.610 1.205 1.780 ;
        RECT 0.605 0.880 0.775 1.610 ;
        RECT 0.575 0.670 0.775 0.880 ;
        RECT 0.605 0.300 0.775 0.670 ;
    END
  END Y
END sky130_as_sc_hs__nor2_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tap_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
        RECT 0.110 1.460 0.340 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.220 0.430 1.020 ;
        RECT 0.090 -0.120 0.400 0.220 ;
      LAYER li1 ;
        RECT 0.120 0.105 0.340 1.000 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__tap_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tieh
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.730 1.840 1.040 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 0.380 1.040 1.630 ;
    END
  END ONE
END sky130_as_sc_hs__tieh

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tiel
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.105 1.040 0.860 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ZERO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 1.140 1.040 2.390 ;
    END
  END ZERO
END sky130_as_sc_hs__tiel
END LIBRARY
