magic
tech sky130A
magscale 1 2
timestamp 1739787816
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 0 22 460 204
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 262 298 292 496
rect 350 298 380 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 262 48 292 178
rect 350 48 380 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 156 166 178
rect 110 72 121 156
rect 155 72 166 156
rect 110 48 166 72
rect 196 150 262 178
rect 196 72 207 150
rect 241 72 262 150
rect 196 48 262 72
rect 292 150 350 178
rect 292 72 303 150
rect 337 72 350 150
rect 292 48 350 72
rect 380 95 433 178
rect 380 61 391 95
rect 425 61 433 95
rect 380 48 433 61
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 298 80 336
rect 110 298 166 496
rect 196 488 262 496
rect 196 406 207 488
rect 241 406 262 488
rect 196 298 262 406
rect 292 474 350 496
rect 292 406 303 474
rect 337 406 350 474
rect 292 298 350 406
rect 380 484 433 496
rect 380 450 391 484
rect 425 450 433 484
rect 380 298 433 450
<< ndiffc >>
rect 35 72 69 150
rect 121 72 155 156
rect 207 72 241 150
rect 303 72 337 150
rect 391 61 425 95
<< pdiffc >>
rect 35 336 69 476
rect 207 406 241 488
rect 303 406 337 474
rect 391 450 425 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 262 496 292 522
rect 350 496 380 522
rect 80 266 110 298
rect 30 250 110 266
rect 30 216 40 250
rect 74 216 110 250
rect 30 200 110 216
rect 80 178 110 200
rect 166 266 196 298
rect 262 266 292 298
rect 350 266 380 298
rect 166 250 220 266
rect 166 216 176 250
rect 210 216 220 250
rect 166 200 220 216
rect 262 250 380 266
rect 262 216 272 250
rect 306 216 380 250
rect 262 200 380 216
rect 166 178 196 200
rect 262 178 292 200
rect 350 178 380 200
rect 80 22 110 48
rect 166 22 196 48
rect 262 22 292 48
rect 350 22 380 48
<< polycont >>
rect 40 216 74 250
rect 176 216 210 250
rect 272 216 306 250
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 35 476 69 492
rect 207 488 241 526
rect 207 390 241 406
rect 303 474 337 490
rect 374 484 442 526
rect 374 450 391 484
rect 425 450 442 484
rect 337 406 400 416
rect 303 390 400 406
rect 312 382 400 390
rect 69 336 289 356
rect 35 322 289 336
rect 35 320 142 322
rect 30 250 74 286
rect 30 216 40 250
rect 30 200 74 216
rect 108 172 142 320
rect 176 250 221 288
rect 210 216 221 250
rect 176 200 221 216
rect 255 266 289 322
rect 255 250 306 266
rect 255 216 272 250
rect 255 200 306 216
rect 35 150 69 166
rect 35 21 69 72
rect 108 156 155 172
rect 340 166 400 382
rect 108 72 121 156
rect 108 56 155 72
rect 207 150 241 166
rect 207 21 241 72
rect 303 154 400 166
rect 303 150 374 154
rect 337 132 374 150
rect 303 56 337 72
rect 374 95 442 98
rect 374 61 391 95
rect 425 61 442 95
rect 374 60 442 61
rect 391 21 425 60
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 B
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__or2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 220
string MASKHINTS_NSDM 0 -38 460 209
string MASKHINTS_PSDM 0 273 460 582
<< end >>
