magic
tech sky130A
magscale 1 2
timestamp 1733848483
<< nwell >>
rect -38 262 314 582
<< pwell >>
rect 0 -18 276 204
<< nmos >>
rect 80 50 110 183
rect 166 50 196 183
<< pmos >>
rect 80 315 110 498
rect 166 315 196 498
<< ndiff >>
rect 27 156 80 183
rect 27 74 35 156
rect 69 74 80 156
rect 27 50 80 74
rect 110 158 166 183
rect 110 76 121 158
rect 155 76 166 158
rect 110 50 166 76
rect 196 168 249 183
rect 196 94 207 168
rect 241 94 249 168
rect 196 50 249 94
<< pdiff >>
rect 27 486 80 498
rect 27 348 35 486
rect 69 348 80 486
rect 27 315 80 348
rect 110 315 166 498
rect 196 476 249 498
rect 196 346 207 476
rect 241 346 249 476
rect 196 315 249 346
<< ndiffc >>
rect 35 74 69 156
rect 121 76 155 158
rect 207 94 241 168
<< pdiffc >>
rect 35 348 69 486
rect 207 346 241 476
<< poly >>
rect 80 498 110 524
rect 166 498 196 524
rect 80 282 110 315
rect 25 266 110 282
rect 25 232 35 266
rect 69 232 110 266
rect 25 216 110 232
rect 80 183 110 216
rect 166 284 196 315
rect 166 268 249 284
rect 166 234 205 268
rect 239 234 249 268
rect 166 218 249 234
rect 166 183 196 218
rect 80 24 110 50
rect 166 24 196 50
<< polycont >>
rect 35 232 69 266
rect 205 234 239 268
<< locali >>
rect 0 561 276 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 526 276 527
rect 35 486 69 526
rect 207 476 241 492
rect 35 322 69 348
rect 121 346 207 356
rect 121 322 241 346
rect 33 266 87 284
rect 33 232 35 266
rect 69 232 87 266
rect 33 216 87 232
rect 121 176 155 322
rect 189 268 241 286
rect 189 234 205 268
rect 239 234 241 268
rect 189 218 241 234
rect 35 156 69 172
rect 115 158 155 176
rect 115 134 121 158
rect 35 21 69 74
rect 121 60 155 76
rect 207 168 241 184
rect 207 21 241 94
rect 0 17 276 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor2_1
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -48 276 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 0 496 276 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 34 238 68 272 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali 204 238 238 272 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 221 255 221 255 0 FreeSans 200 0 0 0 B
flabel locali 119 136 153 170 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel ndiffc 136 153 136 153 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor2_1.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
