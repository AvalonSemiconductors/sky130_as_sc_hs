magic
tech sky130A
magscale 1 2
timestamp 1740408424
<< nwell >>
rect -38 262 774 582
<< pwell >>
rect 0 20 736 204
rect 26 -20 90 20
rect 486 -15 536 20
rect 486 -20 526 -15
<< pmos >>
rect 80 299 110 496
rect 166 299 196 496
rect 252 299 282 496
rect 338 299 368 496
rect 538 299 568 496
rect 624 299 654 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 252 48 282 178
rect 338 48 368 178
rect 538 48 568 178
rect 624 48 654 178
<< ndiff >>
rect 27 166 80 178
rect 27 62 35 166
rect 69 62 80 166
rect 27 48 80 62
rect 110 142 166 178
rect 110 108 121 142
rect 155 108 166 142
rect 110 48 166 108
rect 196 92 252 178
rect 196 58 207 92
rect 241 58 252 92
rect 196 48 252 58
rect 282 132 338 178
rect 282 98 293 132
rect 327 98 338 132
rect 282 48 338 98
rect 368 92 538 178
rect 368 58 380 92
rect 526 58 538 92
rect 368 48 538 58
rect 568 152 624 178
rect 568 118 579 152
rect 613 118 624 152
rect 568 48 624 118
rect 654 166 708 178
rect 654 62 665 166
rect 699 62 708 166
rect 654 48 708 62
<< pdiff >>
rect 27 474 80 496
rect 27 360 35 474
rect 69 360 80 474
rect 27 299 80 360
rect 110 462 166 496
rect 110 428 121 462
rect 155 428 166 462
rect 110 299 166 428
rect 196 474 252 496
rect 196 360 207 474
rect 241 360 252 474
rect 196 299 252 360
rect 282 390 338 496
rect 282 356 293 390
rect 327 356 338 390
rect 282 299 338 356
rect 368 474 430 496
rect 368 440 379 474
rect 413 440 430 474
rect 368 299 430 440
rect 484 422 538 496
rect 484 320 493 422
rect 527 320 538 422
rect 484 299 538 320
rect 568 342 624 496
rect 568 308 579 342
rect 613 308 624 342
rect 568 299 624 308
rect 654 416 708 496
rect 654 314 665 416
rect 699 314 708 416
rect 654 299 708 314
<< ndiffc >>
rect 35 62 69 166
rect 121 108 155 142
rect 207 58 241 92
rect 293 98 327 132
rect 380 58 526 92
rect 579 118 613 152
rect 665 62 699 166
<< pdiffc >>
rect 35 360 69 474
rect 121 428 155 462
rect 207 360 241 474
rect 293 356 327 390
rect 379 440 413 474
rect 493 320 527 422
rect 579 308 613 342
rect 665 314 699 416
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 538 496 568 522
rect 624 496 654 522
rect 80 268 110 299
rect 166 268 196 299
rect 252 268 282 299
rect 338 268 368 299
rect 62 252 196 268
rect 62 218 78 252
rect 170 218 196 252
rect 62 200 196 218
rect 238 252 370 268
rect 538 266 568 299
rect 624 266 654 299
rect 238 218 264 252
rect 358 218 370 252
rect 238 200 370 218
rect 442 252 656 266
rect 442 218 458 252
rect 510 218 656 252
rect 80 178 110 200
rect 166 178 196 200
rect 252 178 282 200
rect 338 178 368 200
rect 442 198 656 218
rect 538 178 568 198
rect 624 178 654 198
rect 80 22 110 48
rect 166 22 196 48
rect 252 22 282 48
rect 338 22 368 48
rect 538 22 568 48
rect 624 22 654 48
<< polycont >>
rect 78 218 170 252
rect 264 218 358 252
rect 458 218 510 252
<< locali >>
rect 0 561 736 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 526 736 527
rect 32 474 72 490
rect 32 360 35 474
rect 69 378 72 474
rect 114 462 162 526
rect 114 428 121 462
rect 155 428 162 462
rect 114 412 162 428
rect 204 474 416 490
rect 204 378 207 474
rect 69 360 207 378
rect 241 456 379 474
rect 241 360 243 456
rect 376 440 379 456
rect 413 440 416 474
rect 376 424 416 440
rect 490 422 704 442
rect 490 390 493 422
rect 32 344 243 360
rect 277 356 293 390
rect 327 356 493 390
rect 62 252 186 268
rect 62 218 78 252
rect 170 218 186 252
rect 248 252 374 268
rect 248 218 264 252
rect 358 218 374 252
rect 422 262 456 322
rect 490 320 493 356
rect 527 416 704 422
rect 527 404 665 416
rect 527 320 530 404
rect 490 302 530 320
rect 574 342 616 358
rect 574 308 579 342
rect 613 308 616 342
rect 574 292 616 308
rect 664 314 665 404
rect 699 314 704 416
rect 664 298 704 314
rect 422 252 526 262
rect 422 218 458 252
rect 510 218 526 252
rect 248 212 374 218
rect 35 166 69 184
rect 574 176 620 292
rect 121 174 620 176
rect 121 152 613 174
rect 121 142 579 152
rect 293 132 327 142
rect 121 92 155 108
rect 207 92 241 108
rect 35 21 69 62
rect 293 82 327 98
rect 380 92 530 108
rect 579 102 613 118
rect 665 166 699 182
rect 207 21 241 58
rect 526 58 530 92
rect 380 21 530 58
rect 665 21 699 62
rect 0 17 736 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 A
flabel locali 255 221 289 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 272 238 272 238 0 FreeSans 200 0 0 0 B
flabel locali 459 221 493 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel polycont 476 238 476 238 0 FreeSans 200 0 0 0 C
flabel locali 578 221 612 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali 595 238 595 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor3_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 736 216
string MASKHINTS_NSDM 0 -38 736 204
string MASKHINTS_PSDM 0 272 736 582
<< end >>
