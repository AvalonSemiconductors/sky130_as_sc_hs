magic
tech sky130A
magscale 1 2
timestamp 1739729467
<< nwell >>
rect -38 262 1050 582
<< pwell >>
rect 22 48 1012 204
rect 26 44 320 48
rect 26 24 90 44
rect 748 24 1012 48
rect 26 22 110 24
rect 808 22 838 24
rect 894 22 924 24
rect 26 -20 90 22
<< pmos >>
rect 80 375 110 496
rect 176 375 206 496
rect 266 375 296 496
rect 416 393 446 496
rect 512 393 542 496
rect 636 339 666 496
rect 722 339 752 496
rect 808 339 838 496
rect 894 339 924 496
<< nmoslvt >>
rect 80 48 110 138
rect 176 48 206 138
rect 266 48 296 138
rect 382 48 412 138
rect 512 48 542 168
rect 636 48 666 178
rect 722 48 752 178
rect 808 48 838 178
rect 894 48 924 178
<< ndiff >>
rect 586 168 636 178
rect 452 138 512 168
rect 27 114 80 138
rect 27 74 35 114
rect 69 74 80 114
rect 27 48 80 74
rect 110 102 176 138
rect 110 64 121 102
rect 155 64 176 102
rect 110 48 176 64
rect 206 48 266 138
rect 296 108 382 138
rect 296 74 308 108
rect 370 74 382 108
rect 296 48 382 74
rect 412 48 512 138
rect 542 92 636 168
rect 542 58 591 92
rect 625 58 636 92
rect 542 48 636 58
rect 666 170 722 178
rect 666 72 677 170
rect 711 72 722 170
rect 666 48 722 72
rect 752 170 808 178
rect 752 62 763 170
rect 797 62 808 170
rect 752 48 808 62
rect 838 170 894 178
rect 838 74 849 170
rect 883 74 894 170
rect 838 48 894 74
rect 924 170 982 178
rect 924 58 935 170
rect 969 58 982 170
rect 924 48 982 58
<< pdiff >>
rect 27 472 80 496
rect 27 410 35 472
rect 69 410 80 472
rect 27 375 80 410
rect 110 488 176 496
rect 110 452 121 488
rect 155 452 176 488
rect 110 375 176 452
rect 206 375 266 496
rect 296 474 416 496
rect 296 418 330 474
rect 382 418 416 474
rect 296 393 416 418
rect 446 393 512 496
rect 542 488 636 496
rect 542 404 574 488
rect 624 404 636 488
rect 542 393 636 404
rect 296 375 349 393
rect 586 339 636 393
rect 666 466 722 496
rect 666 350 677 466
rect 711 350 722 466
rect 666 339 722 350
rect 752 484 808 496
rect 752 388 763 484
rect 797 388 808 484
rect 752 339 808 388
rect 838 476 894 496
rect 838 354 849 476
rect 883 354 894 476
rect 838 339 894 354
rect 924 488 982 496
rect 924 354 935 488
rect 969 354 982 488
rect 924 339 982 354
<< ndiffc >>
rect 35 74 69 114
rect 121 64 155 102
rect 308 74 370 108
rect 591 58 625 92
rect 677 72 711 170
rect 763 62 797 170
rect 849 74 883 170
rect 935 58 969 170
<< pdiffc >>
rect 35 410 69 472
rect 121 452 155 488
rect 330 418 382 474
rect 574 404 624 488
rect 677 350 711 466
rect 763 388 797 484
rect 849 354 883 476
rect 935 354 969 488
<< poly >>
rect 80 496 110 522
rect 176 496 206 522
rect 266 496 296 522
rect 416 496 446 522
rect 512 496 542 522
rect 636 496 666 522
rect 722 496 752 522
rect 808 496 838 522
rect 894 496 924 522
rect 80 228 110 375
rect 176 334 206 375
rect 266 344 296 375
rect 416 362 446 393
rect 416 346 470 362
rect 152 318 206 334
rect 152 284 162 318
rect 196 284 206 318
rect 152 266 206 284
rect 248 328 306 344
rect 248 294 258 328
rect 292 298 306 328
rect 416 312 426 346
rect 460 312 470 346
rect 292 294 374 298
rect 416 296 470 312
rect 248 268 374 294
rect 80 212 134 228
rect 80 178 90 212
rect 124 178 134 212
rect 80 162 134 178
rect 80 138 110 162
rect 176 138 206 266
rect 248 210 302 226
rect 248 176 258 210
rect 292 176 302 210
rect 248 160 302 176
rect 344 194 374 268
rect 512 254 542 393
rect 636 308 666 339
rect 464 244 542 254
rect 464 210 484 244
rect 518 210 542 244
rect 588 302 666 308
rect 722 302 752 339
rect 808 302 838 339
rect 894 302 924 339
rect 588 292 924 302
rect 588 258 598 292
rect 632 258 924 292
rect 588 242 924 258
rect 464 198 542 210
rect 344 164 412 194
rect 512 168 542 198
rect 636 208 924 242
rect 636 178 666 208
rect 722 178 752 208
rect 808 178 838 208
rect 894 178 924 208
rect 266 138 296 160
rect 382 138 412 164
rect 80 22 110 48
rect 176 22 206 48
rect 266 22 296 48
rect 382 22 412 48
rect 512 22 542 48
rect 636 22 666 48
rect 722 22 752 48
rect 808 22 838 48
rect 894 22 924 48
<< polycont >>
rect 162 284 196 318
rect 258 294 292 328
rect 426 312 460 346
rect 90 178 124 212
rect 258 176 292 210
rect 484 210 518 244
rect 598 258 632 292
<< locali >>
rect 0 561 1012 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 526 1012 527
rect 121 488 155 526
rect 22 472 69 488
rect 22 410 35 472
rect 574 488 626 526
rect 121 436 155 452
rect 314 474 398 476
rect 22 402 69 410
rect 314 418 330 474
rect 382 430 398 474
rect 382 418 540 430
rect 22 368 274 402
rect 314 396 540 418
rect 22 132 56 368
rect 240 344 274 368
rect 416 350 470 362
rect 344 346 470 350
rect 90 318 206 334
rect 90 284 162 318
rect 196 284 206 318
rect 90 268 206 284
rect 240 328 292 344
rect 240 294 258 328
rect 240 278 292 294
rect 344 312 426 346
rect 460 312 470 346
rect 506 346 540 396
rect 624 404 626 488
rect 574 388 626 404
rect 677 466 711 486
rect 763 484 797 526
rect 763 372 797 388
rect 849 476 883 492
rect 506 312 630 346
rect 344 296 470 312
rect 572 308 630 312
rect 677 338 711 350
rect 849 338 883 354
rect 935 488 969 526
rect 935 338 969 354
rect 90 226 136 228
rect 90 224 298 226
rect 344 224 384 296
rect 572 292 642 308
rect 90 212 384 224
rect 124 210 384 212
rect 124 178 258 210
rect 90 176 258 178
rect 292 180 384 210
rect 440 244 538 262
rect 440 210 484 244
rect 518 210 538 244
rect 572 258 598 292
rect 632 258 642 292
rect 572 242 642 258
rect 677 248 883 338
rect 292 176 298 180
rect 90 162 298 176
rect 248 160 298 162
rect 440 158 476 210
rect 572 176 606 242
rect 522 142 606 176
rect 677 170 711 248
rect 22 114 69 132
rect 522 124 556 142
rect 22 100 35 114
rect 35 58 69 74
rect 121 102 155 118
rect 121 21 155 64
rect 296 108 556 124
rect 296 74 308 108
rect 370 90 556 108
rect 590 92 628 108
rect 370 74 384 90
rect 296 58 384 74
rect 590 58 591 92
rect 625 58 628 92
rect 590 21 628 58
rect 677 56 711 72
rect 763 170 797 188
rect 763 21 797 62
rect 849 170 883 248
rect 849 58 883 74
rect 935 170 969 192
rect 935 21 969 58
rect 0 17 1012 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 170 170 204 204 0 FreeSans 200 0 0 0 S
port 8 nsew signal input
flabel locali 187 187 187 187 0 FreeSans 200 0 0 0 S
flabel locali 153 289 187 323 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 170 306 170 306 0 FreeSans 200 0 0 0 B
flabel locali 442 221 476 255 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 459 238 459 238 0 FreeSans 200 0 0 0 A
flabel locali 697 255 731 289 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 714 272 714 272 0 FreeSans 200 0 0 0 Y
flabel locali 425 306 459 340 0 FreeSans 200 0 0 0 S
port 8 nsew signal input
flabel locali 442 323 442 323 0 FreeSans 200 0 0 0 S
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__mux2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1012 216
string MASKHINTS_NSDM 0 -34 1012 204
string MASKHINTS_PSDM 0 289 1012 578
<< end >>
