magic
tech sky130A
magscale 1 2
timestamp 1734440952
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 10 48 450 204
rect 26 44 320 48
rect 26 -20 90 44
<< pmos >>
rect 80 316 110 496
rect 166 316 196 496
rect 262 316 292 496
rect 350 316 380 496
<< nmoslvt >>
rect 80 49 110 184
rect 166 49 196 184
rect 262 49 292 184
rect 350 49 380 184
<< ndiff >>
rect 27 168 80 184
rect 27 72 35 168
rect 69 72 80 168
rect 27 49 80 72
rect 110 156 166 184
rect 110 72 121 156
rect 155 72 166 156
rect 110 49 166 72
rect 196 156 262 184
rect 196 72 207 156
rect 241 72 262 156
rect 196 49 262 72
rect 292 168 350 184
rect 292 72 303 168
rect 337 72 350 168
rect 292 49 350 72
rect 380 104 433 184
rect 380 61 391 104
rect 425 61 433 104
rect 380 49 433 61
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 316 80 336
rect 110 316 166 496
rect 196 488 262 496
rect 196 406 207 488
rect 241 406 262 488
rect 196 316 262 406
rect 292 474 350 496
rect 292 406 303 474
rect 337 406 350 474
rect 292 316 350 406
rect 380 484 433 496
rect 380 450 391 484
rect 425 450 433 484
rect 380 316 433 450
<< ndiffc >>
rect 35 72 69 168
rect 121 72 155 156
rect 207 72 241 156
rect 303 72 337 168
rect 391 61 425 104
<< pdiffc >>
rect 35 336 69 476
rect 207 406 241 488
rect 303 406 337 474
rect 391 450 425 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 262 496 292 522
rect 350 496 380 522
rect 80 288 110 316
rect 30 268 110 288
rect 30 234 40 268
rect 74 234 110 268
rect 30 218 110 234
rect 80 184 110 218
rect 166 272 196 316
rect 262 288 292 316
rect 350 288 380 316
rect 166 256 220 272
rect 166 222 176 256
rect 210 222 220 256
rect 166 204 220 222
rect 262 268 380 288
rect 262 234 272 268
rect 306 234 380 268
rect 262 218 380 234
rect 166 184 196 204
rect 262 184 292 218
rect 350 184 380 218
rect 80 23 110 49
rect 166 23 196 49
rect 262 23 292 49
rect 350 23 380 49
<< polycont >>
rect 40 234 74 268
rect 176 222 210 256
rect 272 234 306 268
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 35 476 69 492
rect 207 488 241 526
rect 207 390 241 406
rect 303 474 337 490
rect 374 484 442 526
rect 374 450 391 484
rect 425 450 442 484
rect 337 406 400 416
rect 303 390 400 406
rect 312 382 400 390
rect 69 336 289 356
rect 35 322 289 336
rect 35 320 142 322
rect 30 268 74 286
rect 30 234 40 268
rect 30 218 74 234
rect 35 168 69 184
rect 35 21 69 72
rect 108 172 142 320
rect 255 288 289 322
rect 176 256 221 288
rect 210 222 221 256
rect 176 206 221 222
rect 255 268 306 288
rect 255 234 272 268
rect 255 218 306 234
rect 340 184 400 382
rect 108 156 155 172
rect 108 72 121 156
rect 108 56 155 72
rect 207 156 241 172
rect 207 21 241 72
rect 303 168 400 184
rect 337 154 400 168
rect 337 150 374 154
rect 303 56 337 72
rect 391 104 425 120
rect 391 21 425 61
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 4 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 B
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__or2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
