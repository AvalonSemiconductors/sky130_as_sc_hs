VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__and2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 2.760 1.020 ;
        RECT 0.000 0.110 2.300 0.170 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.760 2.810 ;
        RECT 0.425 1.500 0.595 2.630 ;
        RECT 1.430 2.010 1.600 2.630 ;
        RECT 2.415 1.610 2.585 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.470 0.300 1.810 0.480 ;
        RECT 1.555 0.105 1.725 0.300 ;
        RECT 2.415 0.105 2.585 0.910 ;
        RECT 0.000 -0.085 2.760 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.340 0.990 0.850 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.110 0.990 1.380 1.390 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.480 2.155 2.460 ;
        RECT 1.985 1.070 2.300 1.480 ;
        RECT 1.985 0.600 2.155 1.070 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.880 1.730 1.050 2.250 ;
        RECT 0.880 1.560 1.810 1.730 ;
        RECT 1.640 0.820 1.810 1.560 ;
        RECT 0.355 0.650 1.810 0.820 ;
  END
END sky130_as_sc_hs__and2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__and2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 3.680 1.020 ;
        RECT 0.000 0.110 2.300 0.170 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.425 1.500 0.595 2.630 ;
        RECT 1.430 2.010 1.600 2.630 ;
        RECT 2.415 1.610 2.585 2.630 ;
        RECT 3.280 1.460 3.450 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.470 0.300 1.810 0.480 ;
        RECT 1.555 0.105 1.725 0.300 ;
        RECT 2.415 0.105 2.585 0.910 ;
        RECT 3.300 0.105 3.470 0.930 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.340 0.990 0.850 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.110 0.990 1.380 1.390 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.480 2.155 2.460 ;
        RECT 1.985 1.350 2.300 1.480 ;
        RECT 2.845 1.350 3.015 2.460 ;
        RECT 1.985 1.170 3.015 1.350 ;
        RECT 1.985 1.070 2.300 1.170 ;
        RECT 1.985 0.600 2.155 1.070 ;
        RECT 2.845 0.600 3.015 1.170 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.880 1.730 1.050 2.250 ;
        RECT 0.880 1.560 1.810 1.730 ;
        RECT 1.640 0.820 1.810 1.560 ;
        RECT 0.355 0.650 1.810 0.820 ;
  END
END sky130_as_sc_hs__and2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao21_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 3.220 1.020 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.220 2.810 ;
        RECT 0.605 2.190 0.775 2.630 ;
        RECT 1.985 1.860 2.155 2.630 ;
        RECT 2.845 1.610 3.015 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.280 1.290 0.490 ;
        RECT 1.035 0.105 1.210 0.280 ;
        RECT 1.985 0.105 2.155 0.550 ;
        RECT 2.845 0.105 3.015 0.740 ;
        RECT 0.000 -0.085 3.220 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 0.775 0.440 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.330 0.860 1.680 ;
        RECT 0.610 1.000 1.000 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 1.000 1.510 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.490 2.585 2.460 ;
        RECT 2.415 0.860 2.680 1.490 ;
        RECT 2.415 0.540 2.585 0.860 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.020 0.345 2.370 ;
        RECT 1.035 2.020 1.205 2.370 ;
        RECT 0.175 1.850 1.205 2.020 ;
        RECT 0.175 1.670 0.345 1.850 ;
        RECT 1.035 1.670 1.205 1.850 ;
        RECT 1.465 1.750 1.635 2.290 ;
        RECT 1.465 1.580 1.850 1.750 ;
        RECT 1.680 1.250 1.850 1.580 ;
        RECT 2.050 1.250 2.220 1.330 ;
        RECT 1.680 1.080 2.220 1.250 ;
        RECT 1.680 0.830 1.850 1.080 ;
        RECT 2.050 1.000 2.220 1.080 ;
        RECT 0.610 0.660 1.850 0.830 ;
        RECT 0.175 0.445 0.345 0.605 ;
        RECT 0.610 0.445 0.780 0.660 ;
        RECT 1.465 0.500 1.635 0.660 ;
        RECT 0.175 0.275 0.780 0.445 ;
  END
END sky130_as_sc_hs__ao21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao21_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.140 1.020 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.605 2.190 0.775 2.630 ;
        RECT 1.985 1.860 2.155 2.630 ;
        RECT 2.845 1.610 3.015 2.630 ;
        RECT 3.705 1.470 3.875 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.280 1.290 0.490 ;
        RECT 1.035 0.105 1.210 0.280 ;
        RECT 1.985 0.105 2.155 0.550 ;
        RECT 2.845 0.105 3.015 0.740 ;
        RECT 3.705 0.105 3.875 0.900 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 0.775 0.440 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.330 0.860 1.680 ;
        RECT 0.610 1.000 1.000 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 1.000 1.510 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.490 2.585 2.460 ;
        RECT 2.415 1.310 2.720 1.490 ;
        RECT 3.275 1.310 3.445 2.460 ;
        RECT 2.415 1.090 3.445 1.310 ;
        RECT 2.415 0.860 2.720 1.090 ;
        RECT 2.415 0.280 2.585 0.860 ;
        RECT 3.275 0.290 3.445 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.020 0.345 2.460 ;
        RECT 1.035 2.020 1.205 2.460 ;
        RECT 0.175 1.850 1.205 2.020 ;
        RECT 0.175 1.500 0.345 1.850 ;
        RECT 1.035 1.500 1.205 1.850 ;
        RECT 1.465 1.750 1.635 2.460 ;
        RECT 1.465 1.580 1.850 1.750 ;
        RECT 1.680 1.330 1.850 1.580 ;
        RECT 1.680 1.000 2.240 1.330 ;
        RECT 1.680 0.830 1.850 1.000 ;
        RECT 0.610 0.660 1.850 0.830 ;
        RECT 0.175 0.445 0.345 0.605 ;
        RECT 0.610 0.445 0.780 0.660 ;
        RECT 0.175 0.275 0.780 0.445 ;
        RECT 1.465 0.280 1.635 0.660 ;
  END
END sky130_as_sc_hs__ao21_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao21b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao21b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.130 -0.110 0.340 0.140 ;
        RECT 1.380 0.110 3.680 0.140 ;
        RECT 1.510 -0.100 1.830 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.170 1.500 0.775 2.630 ;
        RECT 1.985 2.190 2.155 2.630 ;
        RECT 3.365 1.860 3.535 2.630 ;
        RECT 4.225 1.610 4.395 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.105 0.775 0.830 ;
        RECT 2.330 0.280 2.670 0.490 ;
        RECT 2.415 0.105 2.590 0.280 ;
        RECT 3.365 0.105 3.535 0.550 ;
        RECT 4.225 0.105 4.395 0.740 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.410 1.000 0.860 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.330 2.240 1.680 ;
        RECT 1.990 1.000 2.380 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.620 1.000 2.890 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 3.795 1.490 3.965 2.460 ;
        RECT 3.795 0.860 4.070 1.490 ;
        RECT 3.795 0.600 3.965 0.860 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.035 1.170 1.205 2.460 ;
        RECT 1.555 2.020 1.725 2.290 ;
        RECT 2.415 2.020 2.585 2.290 ;
        RECT 1.555 1.850 2.585 2.020 ;
        RECT 1.555 1.500 1.725 1.850 ;
        RECT 2.415 1.500 2.585 1.850 ;
        RECT 2.845 1.750 3.015 2.290 ;
        RECT 2.845 1.580 3.230 1.750 ;
        RECT 1.570 1.170 1.820 1.330 ;
        RECT 1.035 1.000 1.820 1.170 ;
        RECT 3.060 1.250 3.230 1.580 ;
        RECT 3.430 1.250 3.600 1.330 ;
        RECT 3.060 1.080 3.600 1.250 ;
        RECT 1.035 0.450 1.205 1.000 ;
        RECT 3.060 0.830 3.230 1.080 ;
        RECT 3.430 1.000 3.600 1.080 ;
        RECT 1.990 0.660 3.230 0.830 ;
        RECT 1.555 0.445 1.725 0.605 ;
        RECT 1.990 0.445 2.160 0.660 ;
        RECT 2.845 0.500 3.015 0.660 ;
        RECT 1.555 0.275 2.160 0.445 ;
  END
END sky130_as_sc_hs__ao21b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao21b_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao21b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 5.520 1.020 ;
        RECT 0.000 0.140 4.600 0.150 ;
        RECT 0.130 -0.110 0.340 0.140 ;
        RECT 1.380 0.110 3.680 0.140 ;
        RECT 1.510 -0.100 1.830 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.520 2.810 ;
        RECT 0.170 1.500 0.775 2.630 ;
        RECT 1.985 2.190 2.155 2.630 ;
        RECT 3.365 1.860 3.535 2.630 ;
        RECT 4.225 1.610 4.395 2.630 ;
        RECT 5.085 1.440 5.255 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.105 0.775 0.830 ;
        RECT 2.330 0.280 2.670 0.450 ;
        RECT 2.415 0.105 2.590 0.280 ;
        RECT 3.365 0.105 3.535 0.550 ;
        RECT 4.225 0.105 4.395 0.740 ;
        RECT 5.085 0.105 5.255 0.930 ;
        RECT 0.000 -0.085 5.520 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.410 1.000 0.860 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.330 2.240 1.680 ;
        RECT 1.990 1.000 2.380 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.620 1.000 2.890 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 3.795 1.490 3.965 2.460 ;
        RECT 3.795 1.250 4.040 1.490 ;
        RECT 4.655 1.250 4.825 2.460 ;
        RECT 3.795 1.040 4.825 1.250 ;
        RECT 3.795 0.860 4.040 1.040 ;
        RECT 3.795 0.600 3.965 0.860 ;
        RECT 4.655 0.600 4.825 1.040 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.035 1.200 1.205 2.260 ;
        RECT 1.555 2.020 1.725 2.290 ;
        RECT 2.415 2.020 2.585 2.290 ;
        RECT 1.555 1.850 2.585 2.020 ;
        RECT 1.555 1.500 1.725 1.850 ;
        RECT 2.415 1.500 2.585 1.850 ;
        RECT 2.845 1.750 3.015 2.290 ;
        RECT 2.845 1.580 3.230 1.750 ;
        RECT 1.570 1.200 1.820 1.330 ;
        RECT 1.035 1.000 1.820 1.200 ;
        RECT 3.060 1.250 3.230 1.580 ;
        RECT 3.430 1.250 3.600 1.330 ;
        RECT 3.060 1.080 3.600 1.250 ;
        RECT 1.035 0.520 1.205 1.000 ;
        RECT 3.060 0.830 3.230 1.080 ;
        RECT 3.430 1.000 3.600 1.080 ;
        RECT 1.990 0.660 3.230 0.830 ;
        RECT 1.555 0.445 1.725 0.605 ;
        RECT 1.990 0.445 2.160 0.660 ;
        RECT 2.845 0.500 3.015 0.660 ;
        RECT 1.555 0.275 2.160 0.445 ;
  END
END sky130_as_sc_hs__ao21b_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao22_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 3.680 1.020 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.605 2.440 0.775 2.630 ;
        RECT 0.520 2.270 0.860 2.440 ;
        RECT 2.475 1.510 2.645 2.630 ;
        RECT 3.335 1.440 3.505 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.960 0.290 1.300 0.480 ;
        RECT 1.045 0.105 1.215 0.290 ;
        RECT 2.475 0.105 2.645 0.830 ;
        RECT 3.335 0.105 3.505 0.930 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 1.340 0.430 1.760 ;
        RECT 0.210 1.000 0.480 1.340 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.160 1.340 1.350 1.760 ;
        RECT 1.160 1.190 1.460 1.340 ;
        RECT 1.240 1.000 1.460 1.190 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.760 1.340 0.990 1.760 ;
        RECT 0.760 1.000 0.980 1.340 ;
    END
  END B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.640 1.000 1.940 1.340 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.490 3.075 2.460 ;
        RECT 2.820 0.920 3.110 1.490 ;
        RECT 2.905 0.280 3.075 0.920 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.100 0.345 2.460 ;
        RECT 1.045 2.290 2.125 2.460 ;
        RECT 1.045 2.100 1.215 2.290 ;
        RECT 1.955 2.130 2.125 2.290 ;
        RECT 0.175 1.930 1.215 2.100 ;
        RECT 1.520 1.830 1.690 2.120 ;
        RECT 1.520 1.660 2.280 1.830 ;
        RECT 2.110 1.340 2.280 1.660 ;
        RECT 2.110 1.000 2.530 1.340 ;
        RECT 2.110 0.830 2.280 1.000 ;
        RECT 0.175 0.660 2.280 0.830 ;
        RECT 0.175 0.280 0.345 0.660 ;
        RECT 1.925 0.300 2.095 0.660 ;
  END
END sky130_as_sc_hs__ao22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao22_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.605 2.440 0.775 2.630 ;
        RECT 0.520 2.270 0.860 2.440 ;
        RECT 2.475 1.510 2.645 2.630 ;
        RECT 3.335 1.440 3.505 2.630 ;
        RECT 4.205 1.440 4.375 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.960 0.290 1.300 0.480 ;
        RECT 1.045 0.105 1.215 0.290 ;
        RECT 2.475 0.105 2.645 0.830 ;
        RECT 3.335 0.105 3.505 0.930 ;
        RECT 4.205 0.105 4.375 0.930 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 1.340 0.430 1.760 ;
        RECT 0.210 1.000 0.480 1.340 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.160 1.340 1.350 1.760 ;
        RECT 1.160 1.190 1.460 1.340 ;
        RECT 1.240 1.000 1.460 1.190 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.760 1.340 0.990 1.760 ;
        RECT 0.760 1.000 0.980 1.340 ;
    END
  END B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.640 1.000 1.940 1.340 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.490 3.075 2.460 ;
        RECT 2.820 1.270 3.110 1.490 ;
        RECT 3.765 1.270 3.935 2.460 ;
        RECT 2.820 1.100 3.935 1.270 ;
        RECT 2.820 0.920 3.110 1.100 ;
        RECT 2.905 0.280 3.075 0.920 ;
        RECT 3.765 0.280 3.935 1.100 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.100 0.345 2.460 ;
        RECT 1.045 2.290 2.125 2.460 ;
        RECT 1.045 2.100 1.215 2.290 ;
        RECT 1.955 2.130 2.125 2.290 ;
        RECT 0.175 1.930 1.215 2.100 ;
        RECT 1.520 1.830 1.690 2.120 ;
        RECT 1.520 1.660 2.280 1.830 ;
        RECT 2.110 1.340 2.280 1.660 ;
        RECT 2.110 1.000 2.530 1.340 ;
        RECT 2.110 0.830 2.280 1.000 ;
        RECT 0.175 0.660 2.280 0.830 ;
        RECT 0.175 0.280 0.345 0.660 ;
        RECT 1.925 0.300 2.095 0.660 ;
  END
END sky130_as_sc_hs__ao22_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao31_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 3.680 1.020 ;
        RECT 0.000 0.140 3.220 0.150 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 1.155 2.440 1.325 2.630 ;
        RECT 1.070 2.260 1.410 2.440 ;
        RECT 2.085 1.510 2.255 2.630 ;
        RECT 3.235 1.620 3.405 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.300 0.425 0.490 ;
        RECT 2.025 0.300 2.365 0.470 ;
        RECT 0.175 0.105 0.345 0.300 ;
        RECT 2.105 0.105 2.275 0.300 ;
        RECT 3.235 0.105 3.405 0.760 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.890 1.000 1.140 1.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.310 1.000 1.670 1.340 ;
        RECT 1.310 0.620 1.510 1.000 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.880 1.000 2.150 1.340 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 1.340 0.710 1.750 ;
        RECT 0.480 1.000 0.710 1.340 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.852800 ;
    PORT
      LAYER li1 ;
        RECT 2.800 1.490 2.970 2.460 ;
        RECT 2.800 0.890 3.120 1.490 ;
        RECT 2.800 0.280 2.970 0.890 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.135 1.490 0.345 2.450 ;
        RECT 0.650 2.090 0.820 2.450 ;
        RECT 1.635 2.090 1.815 2.450 ;
        RECT 0.650 1.920 1.815 2.090 ;
        RECT 0.135 0.830 0.305 1.490 ;
        RECT 2.360 1.000 2.630 1.340 ;
        RECT 0.135 0.660 0.775 0.830 ;
        RECT 2.360 0.810 2.540 1.000 ;
        RECT 0.605 0.450 0.775 0.660 ;
        RECT 1.680 0.640 2.540 0.810 ;
        RECT 1.680 0.450 1.850 0.640 ;
        RECT 0.605 0.280 1.850 0.450 ;
  END
END sky130_as_sc_hs__ao31_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__ao31_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__ao31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 1.155 2.440 1.325 2.630 ;
        RECT 1.070 2.260 1.410 2.440 ;
        RECT 2.085 1.510 2.255 2.630 ;
        RECT 3.235 1.620 3.405 2.630 ;
        RECT 4.095 1.450 4.265 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.300 0.425 0.490 ;
        RECT 2.025 0.300 2.365 0.470 ;
        RECT 0.175 0.105 0.345 0.300 ;
        RECT 2.105 0.105 2.275 0.300 ;
        RECT 3.235 0.105 3.405 0.760 ;
        RECT 4.095 0.105 4.265 0.930 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.890 1.000 1.140 1.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.310 1.000 1.670 1.340 ;
        RECT 1.310 0.620 1.510 1.000 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.880 1.000 2.150 1.340 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 1.340 0.710 1.750 ;
        RECT 0.480 1.000 0.710 1.340 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.312000 ;
    PORT
      LAYER li1 ;
        RECT 2.800 1.490 2.970 2.460 ;
        RECT 2.800 1.300 3.120 1.490 ;
        RECT 3.665 1.300 3.835 2.460 ;
        RECT 2.800 1.080 3.835 1.300 ;
        RECT 2.800 0.890 3.120 1.080 ;
        RECT 2.800 0.280 2.970 0.890 ;
        RECT 3.665 0.280 3.835 1.080 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.135 1.490 0.345 2.450 ;
        RECT 0.650 2.090 0.820 2.450 ;
        RECT 1.635 2.090 1.815 2.450 ;
        RECT 0.650 1.920 1.815 2.090 ;
        RECT 0.135 0.830 0.305 1.490 ;
        RECT 2.360 1.000 2.630 1.340 ;
        RECT 0.135 0.660 0.775 0.830 ;
        RECT 2.360 0.810 2.540 1.000 ;
        RECT 0.605 0.450 0.775 0.660 ;
        RECT 1.680 0.640 2.540 0.810 ;
        RECT 1.680 0.450 1.850 0.640 ;
        RECT 0.605 0.280 1.850 0.450 ;
  END
END sky130_as_sc_hs__ao31_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__aoi211_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__aoi211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.120 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.150 1.500 0.370 2.630 ;
        RECT 1.010 1.960 1.230 2.630 ;
        RECT 1.870 2.170 2.090 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.580 0.105 0.800 0.540 ;
        RECT 2.390 0.105 2.610 0.560 ;
        RECT 3.250 0.105 3.470 0.560 ;
        RECT 4.120 0.105 4.320 0.730 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.490500 ;
    PORT
      LAYER li1 ;
        RECT 1.820 1.280 1.990 1.580 ;
        RECT 1.260 1.080 1.990 1.280 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.424500 ;
    PORT
      LAYER li1 ;
        RECT 2.930 1.280 3.130 1.600 ;
        RECT 2.640 1.080 3.130 1.280 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.424500 ;
    PORT
      LAYER li1 ;
        RECT 4.140 1.330 4.310 1.460 ;
        RECT 3.900 1.080 4.310 1.330 ;
        RECT 4.140 0.900 4.310 1.080 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.695800 ;
    PORT
      LAYER li1 ;
        RECT 3.700 1.670 3.900 2.110 ;
        RECT 3.430 1.500 3.900 1.670 ;
        RECT 3.430 0.910 3.660 1.500 ;
        RECT 1.380 0.730 3.930 0.910 ;
        RECT 1.380 0.680 1.720 0.730 ;
        RECT 2.830 0.280 3.030 0.730 ;
        RECT 2.845 0.275 3.015 0.280 ;
        RECT 3.690 0.275 3.930 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    PORT
      LAYER li1 ;
        RECT 0.550 1.290 0.730 1.440 ;
        RECT 0.170 1.080 0.730 1.290 ;
        RECT 0.550 1.060 0.730 1.080 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.590 1.790 0.790 2.460 ;
        RECT 1.450 1.950 1.650 2.460 ;
        RECT 2.400 2.280 4.320 2.450 ;
        RECT 2.400 2.120 2.600 2.280 ;
        RECT 2.830 1.950 3.040 2.110 ;
        RECT 1.450 1.790 3.040 1.950 ;
        RECT 3.250 1.840 3.470 2.280 ;
        RECT 0.590 1.780 3.040 1.790 ;
        RECT 0.590 1.610 1.650 1.780 ;
        RECT 4.120 1.630 4.320 2.280 ;
        RECT 0.160 0.710 1.210 0.890 ;
        RECT 0.160 0.280 0.370 0.710 ;
        RECT 1.010 0.480 1.210 0.710 ;
        RECT 1.810 0.480 2.150 0.530 ;
        RECT 1.010 0.280 2.150 0.480 ;
  END
END sky130_as_sc_hs__aoi211_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__aoi21_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__aoi21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 3.220 1.020 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.220 2.810 ;
        RECT 0.605 2.100 0.775 2.630 ;
        RECT 1.465 2.100 1.635 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.810 0.280 2.150 0.490 ;
        RECT 1.895 0.105 2.065 0.280 ;
        RECT 2.765 0.105 2.935 0.820 ;
        RECT 0.000 -0.085 3.220 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.380 1.420 1.790 1.590 ;
        RECT 0.380 1.330 0.550 1.420 ;
        RECT 0.300 1.000 0.550 1.330 ;
        RECT 1.620 1.330 1.790 1.420 ;
        RECT 1.620 1.000 1.890 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.830 1.000 1.410 1.250 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.670 0.990 2.920 1.590 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641200 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.580 2.495 2.120 ;
        RECT 2.260 0.830 2.495 1.580 ;
        RECT 1.035 0.660 2.495 0.830 ;
        RECT 1.035 0.280 1.205 0.660 ;
        RECT 2.325 0.280 2.495 0.660 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.930 0.345 2.460 ;
        RECT 1.035 1.930 1.205 2.460 ;
        RECT 1.895 2.290 2.925 2.460 ;
        RECT 1.895 1.930 2.065 2.290 ;
        RECT 0.175 1.760 2.065 1.930 ;
        RECT 2.755 1.760 2.925 2.290 ;
  END
END sky130_as_sc_hs__aoi21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__aoi21b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__aoi21b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 4.140 1.020 ;
        RECT 0.000 0.140 3.220 0.150 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.605 2.100 0.775 2.630 ;
        RECT 1.465 2.100 1.635 2.630 ;
        RECT 3.730 1.500 3.900 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.810 0.280 2.150 0.490 ;
        RECT 1.895 0.105 2.065 0.280 ;
        RECT 2.750 0.105 2.950 0.820 ;
        RECT 3.740 0.105 3.910 0.820 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.380 1.420 1.790 1.590 ;
        RECT 0.380 1.330 0.550 1.420 ;
        RECT 0.300 1.000 0.550 1.330 ;
        RECT 1.620 1.330 1.790 1.420 ;
        RECT 1.620 1.000 1.890 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.830 1.000 1.410 1.250 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.620 0.990 3.830 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641200 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.580 2.495 2.120 ;
        RECT 2.260 0.830 2.495 1.580 ;
        RECT 1.035 0.660 2.495 0.830 ;
        RECT 1.035 0.280 1.205 0.660 ;
        RECT 2.325 0.280 2.495 0.660 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.930 0.345 2.460 ;
        RECT 1.035 1.930 1.205 2.460 ;
        RECT 1.895 2.290 2.925 2.460 ;
        RECT 1.895 1.930 2.065 2.290 ;
        RECT 0.175 1.760 2.065 1.930 ;
        RECT 2.755 1.500 2.925 2.290 ;
        RECT 3.275 1.330 3.445 2.450 ;
        RECT 2.670 0.990 3.445 1.330 ;
        RECT 3.275 0.280 3.445 0.990 ;
  END
END sky130_as_sc_hs__aoi21b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__aoi22_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__aoi22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 2.855 1.890 3.025 2.630 ;
        RECT 3.715 1.890 3.885 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.280 0.855 0.450 ;
        RECT 3.630 0.280 3.970 0.450 ;
        RECT 0.605 0.105 0.775 0.280 ;
        RECT 3.715 0.105 3.885 0.280 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 1.040 0.740 1.300 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.380 1.310 1.690 1.660 ;
        RECT 1.260 1.060 1.780 1.310 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 1.060 3.170 1.310 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.610 1.040 4.300 1.300 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.165900 ;
    PORT
      LAYER li1 ;
        RECT 0.175 1.720 0.345 2.460 ;
        RECT 1.035 1.830 2.065 2.020 ;
        RECT 1.035 1.720 1.205 1.830 ;
        RECT 0.175 1.550 1.205 1.720 ;
        RECT 1.895 1.720 2.065 1.830 ;
        RECT 1.895 1.550 2.190 1.720 ;
        RECT 1.950 0.890 2.190 1.550 ;
        RECT 1.380 0.680 3.110 0.890 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.605 2.290 2.595 2.460 ;
        RECT 0.605 1.890 0.775 2.290 ;
        RECT 1.465 2.190 1.635 2.290 ;
        RECT 2.425 1.720 2.595 2.290 ;
        RECT 3.285 1.720 3.455 2.460 ;
        RECT 4.145 1.720 4.315 2.460 ;
        RECT 2.425 1.550 4.315 1.720 ;
        RECT 0.175 0.620 1.205 0.800 ;
        RECT 0.175 0.280 0.345 0.620 ;
        RECT 1.035 0.450 1.205 0.620 ;
        RECT 3.285 0.700 4.315 0.870 ;
        RECT 1.810 0.450 2.150 0.470 ;
        RECT 1.035 0.280 2.150 0.450 ;
        RECT 2.340 0.450 2.680 0.470 ;
        RECT 3.285 0.450 3.455 0.700 ;
        RECT 4.145 0.540 4.315 0.700 ;
        RECT 2.340 0.280 3.455 0.450 ;
  END
END sky130_as_sc_hs__aoi22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__aoi31_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__aoi31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.605 2.190 0.775 2.630 ;
        RECT 1.465 2.190 1.635 2.630 ;
        RECT 2.885 2.190 3.055 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.300 0.860 0.470 ;
        RECT 3.665 0.300 3.995 0.470 ;
        RECT 0.605 0.105 0.775 0.300 ;
        RECT 3.745 0.105 3.915 0.300 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.270 1.300 0.550 1.600 ;
        RECT 0.270 0.980 0.980 1.300 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 1.330 1.480 1.600 ;
        RECT 1.200 0.980 1.840 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.610 0.990 3.110 1.330 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.280 1.000 3.710 1.360 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.868700 ;
    PORT
      LAYER li1 ;
        RECT 3.745 1.700 3.915 2.120 ;
        RECT 3.745 1.530 4.050 1.700 ;
        RECT 3.880 1.370 4.050 1.530 ;
        RECT 3.880 0.810 4.180 1.370 ;
        RECT 3.315 0.640 4.345 0.810 ;
        RECT 3.315 0.450 3.485 0.640 ;
        RECT 2.330 0.280 3.485 0.450 ;
        RECT 4.175 0.280 4.345 0.640 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.020 0.345 2.460 ;
        RECT 1.035 2.020 1.205 2.460 ;
        RECT 1.895 2.020 2.065 2.460 ;
        RECT 2.455 2.020 2.625 2.460 ;
        RECT 3.315 2.290 4.345 2.460 ;
        RECT 3.315 2.020 3.485 2.290 ;
        RECT 0.175 1.850 3.485 2.020 ;
        RECT 0.175 1.770 0.345 1.850 ;
        RECT 1.035 1.770 1.205 1.850 ;
        RECT 1.895 1.770 2.065 1.850 ;
        RECT 2.455 1.770 2.625 1.850 ;
        RECT 3.315 1.770 3.485 1.850 ;
        RECT 4.175 1.820 4.345 2.290 ;
        RECT 0.175 0.640 1.205 0.810 ;
        RECT 1.385 0.640 3.135 0.810 ;
        RECT 0.175 0.280 0.345 0.640 ;
        RECT 1.035 0.450 1.205 0.640 ;
        RECT 1.035 0.280 2.160 0.450 ;
  END
END sky130_as_sc_hs__aoi31_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_11
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.180 1.890 0.350 2.630 ;
        RECT 1.050 1.955 1.220 2.630 ;
        RECT 1.930 1.960 2.100 2.630 ;
        RECT 2.830 1.810 3.000 2.630 ;
        RECT 3.710 1.810 3.880 2.630 ;
        RECT 4.590 1.810 4.760 2.630 ;
        RECT 5.470 1.810 5.640 2.630 ;
        RECT 6.360 1.810 6.530 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.105 0.350 0.910 ;
        RECT 0.970 0.310 1.300 0.560 ;
        RECT 1.850 0.310 2.180 0.560 ;
        RECT 1.050 0.105 1.220 0.310 ;
        RECT 1.930 0.105 2.100 0.310 ;
        RECT 2.830 0.105 3.000 0.530 ;
        RECT 3.710 0.105 3.880 0.530 ;
        RECT 4.590 0.105 4.760 0.540 ;
        RECT 5.470 0.105 5.640 0.540 ;
        RECT 6.360 0.105 6.530 0.540 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 7.120 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 1.080 1.870 1.445 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.902800 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.640 2.560 2.460 ;
        RECT 3.270 1.640 3.440 2.460 ;
        RECT 4.150 1.640 4.320 2.460 ;
        RECT 5.030 1.640 5.200 2.460 ;
        RECT 5.920 1.640 6.090 2.460 ;
        RECT 6.800 1.795 6.970 2.460 ;
        RECT 6.800 1.640 7.170 1.795 ;
        RECT 2.390 1.470 7.170 1.640 ;
        RECT 6.890 0.880 7.170 1.470 ;
        RECT 2.390 0.810 7.170 0.880 ;
        RECT 2.390 0.710 7.060 0.810 ;
        RECT 2.390 0.440 2.560 0.710 ;
        RECT 3.270 0.450 3.440 0.710 ;
        RECT 4.150 0.500 4.320 0.710 ;
        RECT 5.030 0.390 5.200 0.710 ;
        RECT 5.910 0.500 6.080 0.710 ;
        RECT 6.800 0.500 6.970 0.710 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 2.280 1.030 6.680 1.100 ;
      LAYER li1 ;
        RECT 0.610 1.785 0.780 2.460 ;
        RECT 1.490 1.785 1.660 2.460 ;
        RECT 0.610 1.615 2.220 1.785 ;
        RECT 2.050 1.290 2.220 1.615 ;
        RECT 2.050 1.085 6.720 1.290 ;
        RECT 2.050 0.900 2.220 1.085 ;
        RECT 0.610 0.730 2.220 0.900 ;
        RECT 0.610 0.500 0.780 0.730 ;
        RECT 1.490 0.420 1.660 0.730 ;
  END
END sky130_as_sc_hs__buff_11


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.605 2.050 0.775 2.630 ;
        RECT 1.490 1.630 1.660 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.290 0.860 0.490 ;
        RECT 0.605 0.105 0.775 0.290 ;
        RECT 1.490 0.105 1.660 0.940 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.210 1.810 1.020 ;
        RECT 0.110 0.150 0.450 0.210 ;
        RECT 0.110 0.110 0.550 0.150 ;
        RECT 0.110 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.500 1.480 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.475600 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.980 1.320 2.310 ;
        RECT 1.150 1.490 1.320 1.980 ;
        RECT 1.150 1.230 1.390 1.490 ;
        RECT 1.150 0.690 1.320 1.230 ;
        RECT 1.050 0.360 1.320 0.690 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.880 0.345 2.420 ;
        RECT 0.175 1.710 0.840 1.880 ;
        RECT 0.670 1.370 0.840 1.710 ;
        RECT 0.670 1.000 0.980 1.370 ;
        RECT 0.670 0.830 0.840 1.000 ;
        RECT 0.175 0.660 0.840 0.830 ;
        RECT 0.175 0.450 0.345 0.660 ;
  END
END sky130_as_sc_hs__buff_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.760 2.810 ;
        RECT 0.605 2.050 0.775 2.630 ;
        RECT 1.490 1.690 1.660 2.630 ;
        RECT 2.370 1.690 2.540 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.290 0.860 0.490 ;
        RECT 0.605 0.105 0.775 0.290 ;
        RECT 1.490 0.105 1.660 0.940 ;
        RECT 2.380 0.105 2.550 0.940 ;
        RECT 0.000 -0.085 2.760 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.240 2.720 1.020 ;
        RECT 0.030 0.210 1.810 0.240 ;
        RECT 0.110 0.130 0.450 0.210 ;
        RECT 0.110 0.110 0.550 0.130 ;
        RECT 0.110 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.000 0.420 1.480 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.951200 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.910 1.320 2.240 ;
        RECT 1.150 1.520 1.320 1.910 ;
        RECT 1.930 1.520 2.100 2.450 ;
        RECT 1.150 1.210 2.100 1.520 ;
        RECT 1.150 0.800 1.320 1.210 ;
        RECT 1.050 0.470 1.320 0.800 ;
        RECT 1.930 0.600 2.100 1.210 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.880 0.345 2.420 ;
        RECT 0.175 1.710 0.880 1.880 ;
        RECT 0.710 1.380 0.880 1.710 ;
        RECT 0.710 0.990 0.980 1.380 ;
        RECT 0.710 0.830 0.880 0.990 ;
        RECT 0.175 0.660 0.880 0.830 ;
        RECT 0.175 0.450 0.345 0.660 ;
  END
END sky130_as_sc_hs__buff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_6
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.175 1.670 0.345 2.630 ;
        RECT 1.045 1.650 1.215 2.630 ;
        RECT 1.930 1.950 2.100 2.630 ;
        RECT 2.800 1.630 2.970 2.630 ;
        RECT 3.670 1.630 3.840 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.790 ;
        RECT 1.045 0.105 1.215 0.830 ;
        RECT 1.930 0.105 2.100 0.610 ;
        RECT 2.800 0.105 2.970 0.910 ;
        RECT 3.680 0.105 3.850 0.950 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 4.140 1.020 ;
        RECT 0.110 0.120 0.450 0.130 ;
        RECT 0.110 0.110 0.550 0.120 ;
        RECT 0.110 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.160 0.960 0.430 1.480 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.402200 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.860 1.660 2.460 ;
        RECT 1.490 1.690 1.780 1.860 ;
        RECT 1.610 1.460 1.780 1.690 ;
        RECT 2.370 1.460 2.540 2.450 ;
        RECT 3.230 1.460 3.400 2.450 ;
        RECT 1.610 1.260 3.400 1.460 ;
        RECT 1.610 0.940 1.780 1.260 ;
        RECT 1.590 0.830 1.780 0.940 ;
        RECT 1.490 0.770 1.780 0.830 ;
        RECT 2.370 1.190 3.400 1.260 ;
        RECT 1.490 0.650 1.760 0.770 ;
        RECT 1.490 0.500 1.660 0.650 ;
        RECT 2.370 0.570 2.540 1.190 ;
        RECT 3.230 0.510 3.400 1.190 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.840 0.110 0.990 0.120 ;
        RECT 1.280 0.110 1.430 0.120 ;
        RECT 1.720 0.110 1.870 0.120 ;
        RECT 2.160 0.110 2.310 0.120 ;
        RECT 2.595 0.110 2.745 0.120 ;
        RECT 3.025 0.110 3.175 0.120 ;
        RECT 3.455 0.110 3.605 0.120 ;
      LAYER li1 ;
        RECT 0.600 1.420 0.780 2.460 ;
        RECT 0.600 1.220 1.420 1.420 ;
        RECT 0.600 0.280 0.780 1.220 ;
        RECT 1.190 1.000 1.420 1.220 ;
  END
END sky130_as_sc_hs__buff_6


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_8
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.520 2.810 ;
        RECT 0.175 1.670 0.345 2.630 ;
        RECT 1.045 1.650 1.215 2.630 ;
        RECT 1.930 1.690 2.100 2.630 ;
        RECT 2.800 1.630 2.970 2.630 ;
        RECT 3.670 1.630 3.840 2.630 ;
        RECT 4.565 1.630 4.735 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.790 ;
        RECT 1.045 0.105 1.215 0.960 ;
        RECT 1.930 0.105 2.100 0.610 ;
        RECT 2.800 0.105 2.970 0.910 ;
        RECT 3.680 0.105 3.850 0.950 ;
        RECT 4.565 0.105 4.735 0.950 ;
        RECT 0.000 -0.085 5.520 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 5.520 1.020 ;
        RECT 0.000 0.130 4.140 0.140 ;
        RECT 0.110 0.120 0.450 0.130 ;
        RECT 0.110 0.110 0.550 0.120 ;
        RECT 0.110 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.738000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 0.990 0.430 1.500 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.132000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 1.520 2.540 2.450 ;
        RECT 2.120 1.460 2.540 1.520 ;
        RECT 3.230 1.460 3.400 2.450 ;
        RECT 4.130 1.460 4.300 2.450 ;
        RECT 5.010 1.460 5.210 2.460 ;
        RECT 2.120 1.240 5.210 1.460 ;
        RECT 2.120 1.130 2.540 1.240 ;
        RECT 2.370 0.280 2.540 1.130 ;
        RECT 3.230 0.550 3.400 1.240 ;
        RECT 4.130 1.220 5.210 1.240 ;
        RECT 4.130 0.540 4.300 1.220 ;
        RECT 5.010 0.530 5.210 1.220 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.840 0.110 0.990 0.120 ;
        RECT 1.280 0.110 1.430 0.120 ;
        RECT 1.720 0.110 1.870 0.120 ;
        RECT 2.160 0.110 2.310 0.120 ;
        RECT 2.595 0.110 2.745 0.120 ;
        RECT 3.025 0.110 3.175 0.120 ;
        RECT 3.455 0.110 3.605 0.120 ;
        RECT 3.920 0.110 4.070 0.120 ;
        RECT 4.360 0.110 4.510 0.120 ;
        RECT 4.790 0.110 4.940 0.120 ;
      LAYER li1 ;
        RECT 0.600 1.420 0.780 2.460 ;
        RECT 1.490 1.420 1.660 2.460 ;
        RECT 0.600 1.340 1.660 1.420 ;
        RECT 0.600 1.220 1.890 1.340 ;
        RECT 0.600 0.280 0.780 1.220 ;
        RECT 1.490 1.000 1.890 1.220 ;
        RECT 1.490 0.280 1.660 1.000 ;
  END
END sky130_as_sc_hs__buff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__clkbuff_11
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__clkbuff_11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.130 1.540 0.400 2.630 ;
        RECT 1.000 1.850 1.270 2.630 ;
        RECT 1.880 1.850 2.150 2.630 ;
        RECT 2.780 1.850 3.050 2.630 ;
        RECT 3.660 1.850 3.930 2.630 ;
        RECT 4.540 1.850 4.810 2.630 ;
        RECT 5.420 1.850 5.690 2.630 ;
        RECT 6.310 1.850 6.580 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.105 0.390 0.670 ;
        RECT 1.010 0.105 1.260 0.550 ;
        RECT 1.890 0.105 2.140 0.550 ;
        RECT 2.790 0.105 3.040 0.560 ;
        RECT 3.670 0.105 3.920 0.560 ;
        RECT 4.550 0.105 4.800 0.560 ;
        RECT 5.430 0.105 5.680 0.560 ;
        RECT 6.320 0.105 6.570 0.560 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 7.120 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.855000 ;
    PORT
      LAYER li1 ;
        RECT 0.260 1.070 1.870 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.680 2.610 2.460 ;
        RECT 3.220 1.680 3.490 2.460 ;
        RECT 4.100 1.680 4.370 2.460 ;
        RECT 4.980 1.680 5.250 2.460 ;
        RECT 5.870 1.680 6.140 2.460 ;
        RECT 6.750 1.870 7.020 2.460 ;
        RECT 6.750 1.680 7.200 1.870 ;
        RECT 2.390 1.510 7.200 1.680 ;
        RECT 6.690 0.900 7.200 1.510 ;
        RECT 2.390 0.730 7.200 0.900 ;
        RECT 2.390 0.280 2.600 0.730 ;
        RECT 3.230 0.280 3.480 0.730 ;
        RECT 4.110 0.280 4.360 0.730 ;
        RECT 4.990 0.280 5.240 0.730 ;
        RECT 5.870 0.280 6.120 0.730 ;
        RECT 6.760 0.700 7.200 0.730 ;
        RECT 6.760 0.280 7.010 0.700 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.570 1.680 0.830 2.460 ;
        RECT 1.440 1.680 1.710 2.460 ;
        RECT 0.570 1.510 2.220 1.680 ;
        RECT 2.050 1.340 2.220 1.510 ;
        RECT 2.050 1.070 6.520 1.340 ;
        RECT 2.050 0.900 2.220 1.070 ;
        RECT 0.570 0.720 2.220 0.900 ;
        RECT 0.570 0.280 0.820 0.720 ;
        RECT 1.450 0.280 1.700 0.720 ;
  END
END sky130_as_sc_hs__clkbuff_11


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__clkbuff_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__clkbuff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.760 2.810 ;
        RECT 0.605 2.050 0.775 2.630 ;
        RECT 1.490 1.690 1.660 2.630 ;
        RECT 2.370 1.690 2.540 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.540 ;
        RECT 1.490 0.105 1.660 0.730 ;
        RECT 2.380 0.105 2.550 0.720 ;
        RECT 0.000 -0.085 2.760 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.240 2.720 1.020 ;
        RECT 0.030 0.210 1.810 0.240 ;
        RECT 0.110 -0.100 0.450 0.210 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213750 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.050 0.510 1.540 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.826500 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.910 1.320 2.420 ;
        RECT 1.150 1.520 1.320 1.910 ;
        RECT 1.930 1.520 2.100 2.450 ;
        RECT 1.150 1.130 2.310 1.520 ;
        RECT 1.150 0.800 1.320 1.130 ;
        RECT 1.050 0.290 1.320 0.800 ;
        RECT 1.930 0.280 2.100 1.130 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.880 0.345 2.420 ;
        RECT 0.175 1.710 0.880 1.880 ;
        RECT 0.710 1.350 0.880 1.710 ;
        RECT 0.710 0.970 0.980 1.350 ;
        RECT 0.710 0.880 0.880 0.970 ;
        RECT 0.175 0.710 0.880 0.880 ;
        RECT 0.175 0.290 0.345 0.710 ;
  END
END sky130_as_sc_hs__clkbuff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__clkbuff_8
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__clkbuff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.260 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.070 2.810 ;
        RECT 0.130 1.540 0.400 2.630 ;
        RECT 1.000 1.850 1.270 2.630 ;
        RECT 1.880 1.850 2.150 2.630 ;
        RECT 2.780 1.850 3.050 2.630 ;
        RECT 3.660 1.850 3.930 2.630 ;
        RECT 4.540 1.850 4.810 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.070 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.105 0.390 0.670 ;
        RECT 1.010 0.105 1.260 0.550 ;
        RECT 1.890 0.105 2.140 0.550 ;
        RECT 2.790 0.105 3.040 0.560 ;
        RECT 3.670 0.105 3.920 0.560 ;
        RECT 4.550 0.105 4.800 0.560 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 5.060 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.681500 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.680 1.710 2.460 ;
        RECT 2.390 1.680 2.610 2.460 ;
        RECT 3.220 1.680 3.490 2.460 ;
        RECT 4.100 1.680 4.370 2.460 ;
        RECT 1.490 1.510 4.910 1.680 ;
        RECT 4.050 0.900 4.910 1.510 ;
        RECT 1.490 0.730 4.910 0.900 ;
        RECT 1.490 0.280 1.700 0.730 ;
        RECT 2.390 0.280 2.600 0.730 ;
        RECT 3.230 0.280 3.480 0.730 ;
        RECT 4.110 0.280 4.360 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.427500 ;
    PORT
      LAYER li1 ;
        RECT 0.130 1.070 0.980 1.340 ;
        RECT 0.130 0.840 0.400 1.070 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.570 1.680 0.820 2.460 ;
        RECT 0.570 1.510 1.320 1.680 ;
        RECT 1.150 1.340 1.320 1.510 ;
        RECT 1.150 1.070 3.880 1.340 ;
        RECT 1.150 0.900 1.320 1.070 ;
        RECT 0.570 0.730 1.320 0.900 ;
        RECT 0.570 0.280 0.820 0.730 ;
  END
END sky130_as_sc_hs__clkbuff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.020 7.360 1.020 ;
        RECT 0.120 -0.110 0.520 -0.020 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.360 1.690 6.980 2.630 ;
        RECT 0.600 1.340 0.850 1.690 ;
        RECT 0.560 1.140 0.890 1.340 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 6.390 0.940 6.720 1.520 ;
        RECT 0.360 0.105 6.970 0.940 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_16


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_3
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.020 1.380 1.020 ;
        RECT 0.110 -0.075 0.380 -0.020 ;
        RECT 0.110 -0.110 0.360 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.980 0.580 1.580 ;
        RECT 0.140 0.105 1.210 0.980 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.140 1.830 1.210 2.630 ;
        RECT 0.830 1.150 1.170 1.830 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
END sky130_as_sc_hs__decap_3


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.020 1.840 1.020 ;
        RECT 0.130 -0.100 0.450 -0.020 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.170 1.850 1.670 2.630 ;
        RECT 1.270 1.180 1.610 1.850 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.900 0.580 1.580 ;
        RECT 0.180 0.105 1.660 0.900 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 9.660 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 8.260 0.140 9.660 0.240 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 9.660 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.510 8.515 2.630 ;
        RECT 9.260 1.780 9.430 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.830 ;
        RECT 9.250 0.105 9.420 0.540 ;
        RECT 0.000 -0.085 9.660 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.530 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.457800 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.150 8.110 1.690 ;
        RECT 7.890 0.300 8.110 1.150 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.457800 ;
    PORT
      LAYER li1 ;
        RECT 8.785 1.680 8.955 2.450 ;
        RECT 8.785 1.510 9.120 1.680 ;
        RECT 8.950 1.420 9.120 1.510 ;
        RECT 8.950 1.020 9.230 1.420 ;
        RECT 8.950 0.830 9.120 1.020 ;
        RECT 8.785 0.660 9.120 0.830 ;
        RECT 8.785 0.280 8.955 0.660 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.240 0.610 1.410 1.590 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 1.060 0.280 1.410 0.610 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 7.030 1.350 7.200 2.030 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.330 1.350 ;
        RECT 6.280 1.060 7.330 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 1.030 7.330 1.060 ;
        RECT 7.030 0.790 7.200 1.030 ;
        RECT 8.500 1.000 8.780 1.340 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 1.170 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 1.170 1.590 1.470 1.610 ;
        RECT 0.860 1.020 1.100 1.350 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 0.900 0.630 1.070 1.020 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 7.120 1.020 7.360 1.330 ;
        RECT 8.580 1.020 8.820 1.310 ;
        RECT 7.190 0.850 8.820 1.020 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 0.900 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxbp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxfp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxfp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 8.710 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.740 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 0.000 -0.085 8.740 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.530 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.457800 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.150 8.110 1.690 ;
        RECT 7.890 0.300 8.110 1.150 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.240 0.610 1.410 1.590 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 1.060 0.280 1.410 0.610 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.200 2.030 ;
        RECT 6.280 1.060 7.200 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 0.790 7.200 1.060 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 1.170 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 1.170 1.590 1.470 1.610 ;
        RECT 0.860 1.020 1.100 1.350 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 0.900 0.630 1.070 1.020 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 0.900 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxfp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxfp_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxfp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 9.660 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 8.260 0.140 9.660 0.240 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 9.660 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
        RECT 9.260 1.440 9.430 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 9.230 0.105 9.400 0.950 ;
        RECT 0.000 -0.085 9.660 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.530 ;
    END
  END CLK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.915600 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.300 8.110 1.690 ;
        RECT 8.785 1.300 8.955 2.450 ;
        RECT 7.690 1.150 8.955 1.300 ;
        RECT 7.890 1.080 8.955 1.150 ;
        RECT 7.890 0.300 8.110 1.080 ;
        RECT 8.785 0.280 8.955 1.080 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.240 0.610 1.410 1.590 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 1.060 0.280 1.410 0.610 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.200 2.030 ;
        RECT 6.280 1.060 7.200 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 0.790 7.200 1.060 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 1.170 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 1.170 1.590 1.470 1.610 ;
        RECT 0.860 1.020 1.100 1.350 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 0.900 0.630 1.070 1.020 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 0.900 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxfp_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtn_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 8.710 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.740 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 0.000 -0.085 8.740 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.530 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.457800 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.150 8.110 1.690 ;
        RECT 7.890 0.300 8.110 1.150 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.880 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.880 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 1.240 0.760 1.410 1.750 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.060 0.280 1.410 0.760 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 7.030 1.350 7.200 2.030 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.520 1.350 ;
        RECT 6.280 1.060 7.520 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 1.000 7.520 1.060 ;
        RECT 7.030 0.790 7.200 1.000 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 0.620 1.840 0.860 1.860 ;
        RECT 0.620 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 0.620 1.590 0.970 1.610 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 1.110 0.630 1.340 0.790 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 1.110 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxtn_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtn_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 9.660 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 8.260 0.140 9.660 0.240 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 9.660 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
        RECT 9.260 1.440 9.430 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 9.230 0.105 9.400 0.950 ;
        RECT 0.000 -0.085 9.660 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.530 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.915600 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.300 8.110 1.690 ;
        RECT 8.785 1.300 8.955 2.450 ;
        RECT 7.690 1.150 8.955 1.300 ;
        RECT 7.890 1.080 8.955 1.150 ;
        RECT 7.890 0.300 8.110 1.080 ;
        RECT 8.785 0.280 8.955 1.080 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.880 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.880 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 1.240 0.810 1.410 1.750 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.060 0.280 1.410 0.810 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 7.030 1.350 7.200 2.030 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.520 1.350 ;
        RECT 6.280 1.060 7.520 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 1.000 7.520 1.060 ;
        RECT 7.030 0.790 7.200 1.000 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 0.650 1.840 0.940 1.890 ;
        RECT 0.650 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 0.650 1.560 0.940 1.610 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 1.090 0.630 1.330 0.820 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 1.090 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxtn_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 8.710 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.740 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 0.000 -0.085 8.740 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246750 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.580 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.150 8.110 1.690 ;
        RECT 7.890 0.300 8.110 1.150 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.240 0.610 1.410 1.590 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 1.060 0.280 1.410 0.610 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 7.030 1.350 7.200 2.030 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.520 1.350 ;
        RECT 6.280 1.060 7.520 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 1.000 7.520 1.060 ;
        RECT 7.030 0.790 7.200 1.000 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 2.410 1.840 2.660 1.880 ;
        RECT 1.170 1.670 4.390 1.840 ;
        RECT 1.170 1.590 1.470 1.670 ;
        RECT 2.410 1.640 2.660 1.670 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.470 1.670 ;
        RECT 4.210 1.320 4.390 1.670 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 0.550 0.630 0.920 0.840 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 0.550 0.580 6.000 0.630 ;
        RECT 0.750 0.490 6.000 0.580 ;
  END
END sky130_as_sc_hs__dfxtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 9.660 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 8.260 0.140 9.660 0.240 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 9.660 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.470 8.515 2.630 ;
        RECT 9.260 1.440 9.430 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.280 0.870 0.470 ;
        RECT 0.620 0.105 0.790 0.280 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.830 ;
        RECT 8.345 0.105 8.515 0.910 ;
        RECT 9.230 0.105 9.400 0.950 ;
        RECT 0.000 -0.085 9.660 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246750 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.980 0.440 1.580 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.300 8.110 1.690 ;
        RECT 8.785 1.300 8.955 2.450 ;
        RECT 7.690 1.150 8.955 1.300 ;
        RECT 7.890 1.080 8.955 1.150 ;
        RECT 7.890 0.300 8.110 1.080 ;
        RECT 8.785 0.280 8.955 1.080 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.161250 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.880 1.680 ;
    END
  END D
  OBS
      LAYER pwell ;
        RECT 8.580 0.110 8.730 0.120 ;
        RECT 9.010 0.110 9.160 0.120 ;
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 2.080 2.070 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.350 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.020 1.070 1.350 ;
        RECT 0.610 0.810 0.780 1.020 ;
        RECT 0.190 0.640 0.780 0.810 ;
        RECT 0.190 0.280 0.360 0.640 ;
        RECT 1.240 0.610 1.410 1.590 ;
        RECT 2.050 1.720 2.250 2.070 ;
        RECT 2.050 0.880 2.220 1.720 ;
        RECT 2.420 1.520 2.630 1.850 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.810 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.390 0.990 2.600 1.320 ;
        RECT 2.050 0.690 2.250 0.880 ;
        RECT 2.800 0.820 2.970 1.610 ;
        RECT 4.170 1.480 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.440 5.100 1.830 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 1.060 0.280 1.410 0.610 ;
        RECT 2.080 0.280 2.250 0.690 ;
        RECT 2.710 0.650 2.970 0.820 ;
        RECT 2.710 0.600 2.880 0.650 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 0.940 5.110 1.270 ;
        RECT 5.280 0.650 5.450 1.620 ;
        RECT 6.670 1.410 6.860 1.620 ;
        RECT 7.030 1.350 7.200 2.030 ;
        RECT 5.790 0.880 6.000 1.240 ;
        RECT 6.280 1.230 6.490 1.240 ;
        RECT 7.030 1.230 7.520 1.350 ;
        RECT 6.280 1.060 7.520 1.230 ;
        RECT 6.280 0.900 6.490 1.060 ;
        RECT 7.030 1.000 7.520 1.060 ;
        RECT 7.030 0.790 7.200 1.000 ;
        RECT 5.190 0.600 5.450 0.650 ;
        RECT 5.030 0.430 5.450 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 2.410 1.840 2.660 1.870 ;
        RECT 1.170 1.670 4.390 1.840 ;
        RECT 1.170 1.590 1.470 1.670 ;
        RECT 2.410 1.640 2.660 1.670 ;
        RECT 2.370 1.100 2.660 1.340 ;
        RECT 3.300 1.190 3.520 1.670 ;
        RECT 4.210 1.320 4.390 1.670 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.660 1.100 ;
        RECT 0.540 0.630 0.840 0.840 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.030 5.170 1.150 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.500 0.630 6.000 0.640 ;
        RECT 0.540 0.610 6.000 0.630 ;
        RECT 0.620 0.490 6.000 0.610 ;
  END
END sky130_as_sc_hs__dfxtp_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__diode_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.220 0.870 1.020 ;
        RECT 0.210 -0.075 0.390 0.220 ;
    END
  END VNB
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.406350 ;
    PORT
      LAYER li1 ;
        RECT 0.190 0.290 0.740 2.450 ;
    END
  END DIODE
END sky130_as_sc_hs__diode_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dyn_dfxtn_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dyn_dfxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 7.820 1.020 ;
        RECT 0.000 0.120 5.520 0.170 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.820 2.810 ;
        RECT 0.660 1.840 0.830 2.630 ;
        RECT 2.365 1.840 2.535 2.630 ;
        RECT 4.515 1.830 4.685 2.630 ;
        RECT 6.495 1.470 6.665 2.630 ;
        RECT 7.355 1.780 7.525 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.320 0.900 0.490 ;
        RECT 2.280 0.320 2.620 0.490 ;
        RECT 4.430 0.320 4.770 0.490 ;
        RECT 6.410 0.320 6.750 0.490 ;
        RECT 0.650 0.105 0.820 0.320 ;
        RECT 2.365 0.105 2.535 0.320 ;
        RECT 4.515 0.105 4.685 0.320 ;
        RECT 6.495 0.105 6.665 0.320 ;
        RECT 7.355 0.105 7.525 0.930 ;
        RECT 0.000 -0.085 7.820 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 1.000 0.770 1.330 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220500 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.000 2.490 1.330 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 6.925 1.590 7.095 2.460 ;
        RECT 6.925 1.100 7.420 1.590 ;
        RECT 6.925 0.580 7.095 1.100 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.175 0.830 0.345 2.460 ;
        RECT 1.000 0.830 1.170 1.970 ;
        RECT 0.175 0.660 1.170 0.830 ;
        RECT 0.175 0.580 0.345 0.660 ;
        RECT 1.340 0.580 1.510 2.460 ;
        RECT 1.865 0.830 2.035 2.460 ;
        RECT 3.990 1.340 4.160 2.460 ;
        RECT 2.690 0.830 2.860 1.330 ;
        RECT 3.170 0.990 3.340 1.330 ;
        RECT 3.650 0.990 3.820 1.330 ;
        RECT 3.990 1.000 4.300 1.340 ;
        RECT 5.970 1.330 6.140 2.460 ;
        RECT 1.865 0.660 2.860 0.830 ;
        RECT 1.865 0.410 2.035 0.660 ;
        RECT 3.990 0.580 4.160 1.000 ;
        RECT 5.150 0.990 5.320 1.330 ;
        RECT 5.630 0.990 5.800 1.330 ;
        RECT 5.970 0.990 6.280 1.330 ;
        RECT 5.970 0.580 6.140 0.990 ;
      LAYER met1 ;
        RECT 1.150 2.000 3.340 2.040 ;
        RECT 0.940 1.870 3.340 2.000 ;
        RECT 0.940 1.770 1.290 1.870 ;
        RECT 3.170 1.750 3.340 1.870 ;
        RECT 3.170 1.580 5.800 1.750 ;
        RECT 3.170 1.330 3.340 1.580 ;
        RECT 5.630 1.330 5.800 1.580 ;
        RECT 3.140 1.020 3.370 1.330 ;
        RECT 3.620 1.020 3.850 1.310 ;
        RECT 5.100 1.030 5.370 1.310 ;
        RECT 1.300 0.550 1.550 0.890 ;
        RECT 3.650 0.550 3.820 1.020 ;
        RECT 5.150 0.550 5.320 1.030 ;
        RECT 5.580 1.020 5.850 1.330 ;
        RECT 1.340 0.380 5.320 0.550 ;
  END
END sky130_as_sc_hs__dyn_dfxtn_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dyn_dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dyn_dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 7.820 1.020 ;
        RECT 0.000 0.120 5.520 0.170 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.820 2.810 ;
        RECT 0.660 1.840 0.830 2.630 ;
        RECT 2.365 1.840 2.535 2.630 ;
        RECT 4.515 1.830 4.685 2.630 ;
        RECT 6.495 1.470 6.665 2.630 ;
        RECT 7.355 1.780 7.525 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.320 0.900 0.490 ;
        RECT 2.280 0.320 2.620 0.490 ;
        RECT 4.430 0.320 4.770 0.490 ;
        RECT 6.410 0.320 6.750 0.490 ;
        RECT 0.650 0.105 0.820 0.320 ;
        RECT 2.365 0.105 2.535 0.320 ;
        RECT 4.515 0.105 4.685 0.320 ;
        RECT 6.495 0.105 6.665 0.320 ;
        RECT 7.355 0.105 7.525 0.930 ;
        RECT 0.000 -0.085 7.820 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 1.000 0.770 1.330 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220500 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.000 2.490 1.330 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 6.925 1.590 7.095 2.460 ;
        RECT 6.925 1.100 7.420 1.590 ;
        RECT 6.925 0.580 7.095 1.100 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.175 0.830 0.345 2.460 ;
        RECT 1.000 0.830 1.170 1.330 ;
        RECT 0.175 0.660 1.170 0.830 ;
        RECT 0.175 0.580 0.345 0.660 ;
        RECT 1.340 0.580 1.510 2.460 ;
        RECT 1.865 0.830 2.035 2.460 ;
        RECT 3.990 1.340 4.160 2.460 ;
        RECT 2.690 0.830 2.860 1.330 ;
        RECT 3.170 0.990 3.340 1.330 ;
        RECT 3.650 0.990 3.820 1.330 ;
        RECT 3.990 1.000 4.300 1.340 ;
        RECT 5.970 1.330 6.140 2.460 ;
        RECT 1.865 0.660 2.860 0.830 ;
        RECT 1.865 0.410 2.035 0.660 ;
        RECT 3.990 0.580 4.160 1.000 ;
        RECT 5.150 0.990 5.320 1.330 ;
        RECT 5.630 0.990 5.800 1.330 ;
        RECT 5.970 0.990 6.280 1.330 ;
        RECT 5.970 0.580 6.140 0.990 ;
      LAYER met1 ;
        RECT 1.280 2.040 1.540 2.080 ;
        RECT 1.280 1.870 3.340 2.040 ;
        RECT 1.280 1.830 1.540 1.870 ;
        RECT 3.170 1.750 3.340 1.870 ;
        RECT 3.170 1.580 5.800 1.750 ;
        RECT 3.170 1.330 3.340 1.580 ;
        RECT 5.630 1.330 5.800 1.580 ;
        RECT 3.140 1.020 3.370 1.330 ;
        RECT 3.620 1.020 3.850 1.310 ;
        RECT 5.100 1.030 5.370 1.310 ;
        RECT 0.970 0.550 1.200 0.890 ;
        RECT 3.650 0.550 3.820 1.020 ;
        RECT 5.150 0.550 5.320 1.030 ;
        RECT 5.580 1.020 5.850 1.330 ;
        RECT 0.970 0.380 5.320 0.550 ;
  END
END sky130_as_sc_hs__dyn_dfxtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dyn_dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dyn_dfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 8.740 1.020 ;
        RECT 0.000 0.120 5.520 0.170 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.740 2.810 ;
        RECT 0.660 1.840 0.830 2.630 ;
        RECT 2.365 1.840 2.535 2.630 ;
        RECT 4.515 1.830 4.685 2.630 ;
        RECT 6.495 1.430 6.665 2.630 ;
        RECT 7.355 1.780 7.525 2.630 ;
        RECT 8.215 1.460 8.385 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.320 0.900 0.490 ;
        RECT 2.280 0.320 2.620 0.490 ;
        RECT 4.430 0.320 4.770 0.490 ;
        RECT 6.410 0.320 6.750 0.490 ;
        RECT 0.650 0.105 0.820 0.320 ;
        RECT 2.365 0.105 2.535 0.320 ;
        RECT 4.515 0.105 4.685 0.320 ;
        RECT 6.495 0.105 6.665 0.320 ;
        RECT 7.355 0.105 7.525 0.930 ;
        RECT 8.215 0.105 8.385 0.930 ;
        RECT 0.000 -0.085 8.740 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 1.000 0.770 1.330 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.220500 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.000 2.490 1.330 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 6.925 1.590 7.095 2.460 ;
        RECT 6.925 1.420 7.420 1.590 ;
        RECT 7.785 1.420 7.955 2.460 ;
        RECT 6.925 1.230 7.955 1.420 ;
        RECT 6.925 1.100 7.420 1.230 ;
        RECT 6.925 0.580 7.095 1.100 ;
        RECT 7.785 0.580 7.955 1.230 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.175 0.830 0.345 2.460 ;
        RECT 1.000 0.830 1.170 1.330 ;
        RECT 0.175 0.660 1.170 0.830 ;
        RECT 0.175 0.580 0.345 0.660 ;
        RECT 1.340 0.580 1.510 2.460 ;
        RECT 1.865 0.830 2.035 2.460 ;
        RECT 3.990 1.340 4.160 2.460 ;
        RECT 2.690 0.830 2.860 1.330 ;
        RECT 3.170 0.990 3.340 1.330 ;
        RECT 3.650 0.990 3.820 1.330 ;
        RECT 3.990 1.000 4.300 1.340 ;
        RECT 5.970 1.330 6.140 2.460 ;
        RECT 1.865 0.660 2.860 0.830 ;
        RECT 1.865 0.410 2.035 0.660 ;
        RECT 3.990 0.580 4.160 1.000 ;
        RECT 5.150 0.990 5.320 1.330 ;
        RECT 5.630 0.990 5.800 1.330 ;
        RECT 5.970 0.990 6.280 1.330 ;
        RECT 5.970 0.580 6.140 0.990 ;
      LAYER met1 ;
        RECT 1.280 2.040 1.540 2.080 ;
        RECT 1.280 1.870 3.340 2.040 ;
        RECT 1.280 1.830 1.540 1.870 ;
        RECT 3.170 1.750 3.340 1.870 ;
        RECT 3.170 1.580 5.800 1.750 ;
        RECT 3.170 1.330 3.340 1.580 ;
        RECT 5.630 1.330 5.800 1.580 ;
        RECT 3.140 1.020 3.370 1.330 ;
        RECT 3.620 1.020 3.850 1.310 ;
        RECT 5.100 1.030 5.370 1.310 ;
        RECT 0.970 0.550 1.200 0.890 ;
        RECT 3.650 0.550 3.820 1.020 ;
        RECT 5.150 0.550 5.320 1.030 ;
        RECT 5.580 1.020 5.850 1.330 ;
        RECT 0.970 0.380 5.320 0.550 ;
  END
END sky130_as_sc_hs__dyn_dfxtp_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_1


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.730 2.020 0.970 2.260 ;
        RECT 0.490 1.780 1.210 2.020 ;
        RECT 0.490 1.300 0.730 1.780 ;
        RECT 0.970 1.300 1.210 1.780 ;
        RECT 1.690 1.540 1.930 2.260 ;
        RECT 3.130 1.540 3.370 2.260 ;
        RECT 4.090 2.020 4.330 2.260 ;
        RECT 1.690 1.300 2.170 1.540 ;
        RECT 0.490 1.060 1.210 1.300 ;
        RECT 0.250 0.820 0.730 1.060 ;
        RECT 0.970 0.820 1.450 1.060 ;
        RECT 0.250 0.340 0.490 0.820 ;
        RECT 1.210 0.340 1.450 0.820 ;
        RECT 1.930 0.820 2.170 1.300 ;
        RECT 2.410 0.820 2.650 1.540 ;
        RECT 2.890 1.300 3.370 1.540 ;
        RECT 3.850 1.780 4.570 2.020 ;
        RECT 3.850 1.300 4.090 1.780 ;
        RECT 4.330 1.300 4.570 1.780 ;
        RECT 5.050 1.540 5.290 2.260 ;
        RECT 6.490 1.540 6.730 2.260 ;
        RECT 5.050 1.300 5.530 1.540 ;
        RECT 2.890 0.820 3.130 1.300 ;
        RECT 3.850 1.060 4.570 1.300 ;
        RECT 1.930 0.580 3.130 0.820 ;
        RECT 3.610 0.820 4.090 1.060 ;
        RECT 4.330 0.820 4.810 1.060 ;
        RECT 2.170 0.340 2.410 0.580 ;
        RECT 2.650 0.340 2.890 0.580 ;
        RECT 3.610 0.340 3.850 0.820 ;
        RECT 4.570 0.340 4.810 0.820 ;
        RECT 5.290 0.820 5.530 1.300 ;
        RECT 5.770 0.820 6.010 1.540 ;
        RECT 6.250 1.300 6.730 1.540 ;
        RECT 6.250 0.820 6.490 1.300 ;
        RECT 5.290 0.580 6.490 0.820 ;
        RECT 5.530 0.340 5.770 0.580 ;
        RECT 6.010 0.340 6.250 0.580 ;
  END
END sky130_as_sc_hs__fill_16


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__hcf_10
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__hcf_10 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.160 5.060 1.020 ;
        RECT 0.000 0.140 4.600 0.160 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.060 2.810 ;
        RECT 0.605 0.280 0.775 2.630 ;
        RECT 1.465 0.280 1.635 2.630 ;
        RECT 2.325 0.290 2.495 2.630 ;
        RECT 3.185 0.290 3.355 2.630 ;
        RECT 4.045 0.290 4.215 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.940 ;
        RECT 1.035 0.105 1.205 0.940 ;
        RECT 1.895 0.105 2.065 0.930 ;
        RECT 2.755 0.105 2.925 0.930 ;
        RECT 3.615 0.105 3.785 0.930 ;
        RECT 4.475 0.105 4.645 0.930 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN HCF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.975000 ;
    PORT
      LAYER li1 ;
        RECT 0.160 1.110 0.435 1.940 ;
    END
  END HCF
END sky130_as_sc_hs__hcf_10


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__iao211_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__iao211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 5.060 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 3.750 0.110 3.900 0.140 ;
        RECT 4.180 0.110 4.330 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.060 2.810 ;
        RECT 0.605 2.080 0.775 2.630 ;
        RECT 2.550 2.190 2.720 2.630 ;
        RECT 3.525 1.850 3.695 2.630 ;
        RECT 4.460 1.580 4.630 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.890 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.895 0.105 2.065 0.540 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.060 0.710 1.300 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.640 1.280 1.870 1.580 ;
        RECT 1.260 1.060 1.870 1.280 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.610 1.320 2.840 1.580 ;
        RECT 2.610 1.060 3.220 1.320 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 4.460 1.300 4.660 1.410 ;
        RECT 4.270 1.060 4.660 1.300 ;
        RECT 4.460 0.850 4.660 1.060 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.013600 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.920 1.635 2.080 ;
        RECT 3.095 1.920 3.265 2.250 ;
        RECT 1.465 1.750 3.265 1.920 ;
        RECT 3.095 1.660 3.265 1.750 ;
        RECT 3.955 1.660 4.125 2.460 ;
        RECT 3.095 1.490 4.125 1.660 ;
        RECT 3.870 1.450 4.125 1.490 ;
        RECT 3.870 0.870 4.090 1.450 ;
        RECT 3.870 0.680 4.210 0.870 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.910 0.345 2.460 ;
        RECT 1.035 2.280 2.065 2.460 ;
        RECT 1.035 1.910 1.205 2.280 ;
        RECT 1.895 2.090 2.065 2.280 ;
        RECT 0.175 1.740 1.205 1.910 ;
        RECT 0.605 0.720 2.410 0.890 ;
        RECT 0.605 0.560 0.775 0.720 ;
        RECT 1.465 0.560 1.635 0.720 ;
        RECT 2.240 0.480 2.410 0.720 ;
        RECT 2.580 0.720 3.695 0.890 ;
        RECT 2.580 0.680 2.915 0.720 ;
        RECT 3.095 0.480 3.265 0.550 ;
        RECT 2.240 0.470 3.265 0.480 ;
        RECT 3.525 0.470 3.695 0.720 ;
        RECT 4.420 0.470 4.590 0.630 ;
        RECT 2.240 0.310 3.350 0.470 ;
        RECT 3.000 0.300 3.350 0.310 ;
        RECT 3.525 0.300 4.590 0.470 ;
  END
END sky130_as_sc_hs__iao211_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 1.380 1.020 ;
        RECT 0.130 -0.075 0.380 0.110 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.030 0.105 1.210 0.940 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.175 1.720 0.345 2.630 ;
        RECT 1.030 1.450 1.210 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.410 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.400 0.775 2.460 ;
        RECT 0.580 0.940 0.790 1.400 ;
        RECT 0.605 0.530 0.775 0.940 ;
    END
  END Y
END sky130_as_sc_hs__inv_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 2.300 1.020 ;
        RECT 0.130 -0.075 0.380 0.110 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.035 0.105 1.205 0.940 ;
        RECT 1.940 0.105 2.110 0.940 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 0.175 1.510 0.345 2.630 ;
        RECT 1.035 1.510 1.205 2.630 ;
        RECT 1.940 1.510 2.110 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.410 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.951200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.340 0.775 2.460 ;
        RECT 0.590 1.310 0.790 1.340 ;
        RECT 1.475 1.310 1.645 2.460 ;
        RECT 0.590 1.110 1.645 1.310 ;
        RECT 0.590 1.000 0.790 1.110 ;
        RECT 0.605 0.530 0.775 1.000 ;
        RECT 1.475 0.520 1.645 1.110 ;
    END
  END Y
END sky130_as_sc_hs__inv_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_6
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 3.220 1.020 ;
        RECT 0.000 0.120 2.300 0.130 ;
        RECT 0.000 0.110 2.320 0.120 ;
        RECT 0.130 -0.075 0.380 0.110 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.410 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.035 0.105 1.205 0.940 ;
        RECT 1.940 0.105 2.110 0.940 ;
        RECT 2.835 0.105 3.005 0.940 ;
        RECT 0.000 -0.085 3.220 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.220 2.810 ;
        RECT 0.175 1.510 0.345 2.630 ;
        RECT 1.035 1.510 1.205 2.630 ;
        RECT 1.940 1.510 2.110 2.630 ;
        RECT 2.825 1.410 2.995 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.476000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.410 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.443200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.340 0.775 2.460 ;
        RECT 0.590 1.310 0.775 1.340 ;
        RECT 1.475 1.310 1.645 2.460 ;
        RECT 2.385 1.310 2.555 2.460 ;
        RECT 0.590 1.110 2.555 1.310 ;
        RECT 0.590 1.000 0.775 1.110 ;
        RECT 0.605 0.600 0.775 1.000 ;
        RECT 1.475 0.600 1.645 1.110 ;
        RECT 2.385 0.600 2.555 1.110 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 2.620 0.110 2.770 0.120 ;
  END
END sky130_as_sc_hs__inv_6


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__maj3_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.140 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.965 2.190 1.135 2.630 ;
        RECT 2.545 2.190 2.715 2.630 ;
        RECT 3.720 1.450 3.890 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.105 1.135 0.540 ;
        RECT 2.600 0.105 2.770 0.540 ;
        RECT 3.720 0.105 3.890 0.900 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.760 1.070 1.280 1.330 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.350 1.500 2.510 1.670 ;
        RECT 0.350 1.330 0.550 1.500 ;
        RECT 0.220 1.070 0.550 1.330 ;
        RECT 2.340 1.330 2.510 1.500 ;
        RECT 2.340 1.070 2.670 1.330 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.550 1.070 2.130 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 3.085 2.240 3.255 2.400 ;
        RECT 3.085 2.070 3.550 2.240 ;
        RECT 3.380 1.310 3.550 2.070 ;
        RECT 3.380 1.040 3.620 1.310 ;
        RECT 3.380 0.550 3.550 1.040 ;
        RECT 3.000 0.380 3.550 0.550 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.170 2.020 0.350 2.300 ;
        RECT 1.750 2.020 1.930 2.460 ;
        RECT 0.170 1.860 2.850 2.020 ;
        RECT 0.170 1.850 3.010 1.860 ;
        RECT 2.680 1.690 3.010 1.850 ;
        RECT 2.840 1.330 3.010 1.690 ;
        RECT 2.840 1.070 3.210 1.330 ;
        RECT 2.840 0.900 3.010 1.070 ;
        RECT 0.175 0.720 3.010 0.900 ;
        RECT 0.175 0.450 0.345 0.720 ;
        RECT 1.755 0.600 1.925 0.720 ;
  END
END sky130_as_sc_hs__maj3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__maj3_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__maj3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 5.060 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.060 2.810 ;
        RECT 0.965 2.190 1.135 2.630 ;
        RECT 2.545 2.190 2.715 2.630 ;
        RECT 3.720 1.470 3.890 2.630 ;
        RECT 4.630 1.450 4.800 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.105 1.135 0.540 ;
        RECT 2.600 0.105 2.770 0.540 ;
        RECT 3.720 0.105 3.890 0.890 ;
        RECT 4.640 0.105 4.810 0.930 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.760 1.070 1.270 1.330 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.500 2.510 1.670 ;
        RECT 0.360 1.330 0.550 1.500 ;
        RECT 0.220 1.070 0.550 1.330 ;
        RECT 2.340 1.330 2.510 1.500 ;
        RECT 2.340 1.070 2.670 1.330 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.550 1.070 2.110 1.330 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 3.085 2.080 3.255 2.280 ;
        RECT 3.085 1.910 3.550 2.080 ;
        RECT 3.380 1.300 3.550 1.910 ;
        RECT 4.155 1.300 4.325 2.450 ;
        RECT 3.380 1.090 4.325 1.300 ;
        RECT 3.380 0.550 3.550 1.090 ;
        RECT 3.000 0.380 3.550 0.550 ;
        RECT 4.155 0.490 4.325 1.090 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 3.950 0.110 4.100 0.120 ;
        RECT 4.380 0.110 4.530 0.120 ;
      LAYER li1 ;
        RECT 0.170 2.020 0.350 2.180 ;
        RECT 1.750 2.020 1.930 2.460 ;
        RECT 0.170 1.850 2.850 2.020 ;
        RECT 2.680 1.750 2.850 1.850 ;
        RECT 2.680 1.500 3.010 1.750 ;
        RECT 2.840 1.330 3.010 1.500 ;
        RECT 2.840 1.000 3.130 1.330 ;
        RECT 2.840 0.900 3.010 1.000 ;
        RECT 0.175 0.730 3.010 0.900 ;
        RECT 0.175 0.470 0.345 0.730 ;
        RECT 1.755 0.600 1.925 0.730 ;
  END
END sky130_as_sc_hs__maj3_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__mux2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.160 4.600 1.020 ;
        RECT 0.000 0.120 4.590 0.160 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.780 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.650 2.170 0.820 2.630 ;
        RECT 3.095 2.170 3.265 2.630 ;
        RECT 4.115 1.570 4.285 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.280 0.860 0.450 ;
        RECT 3.060 0.300 3.400 0.470 ;
        RECT 0.595 0.105 0.775 0.280 ;
        RECT 3.130 0.105 3.310 0.300 ;
        RECT 4.115 0.105 4.285 0.920 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 1.330 2.580 1.640 ;
        RECT 0.450 0.990 0.720 1.330 ;
        RECT 0.550 0.820 0.720 0.990 ;
        RECT 1.420 0.820 1.590 1.330 ;
        RECT 2.330 0.990 2.590 1.330 ;
        RECT 2.380 0.820 2.550 0.990 ;
        RECT 0.550 0.650 2.550 0.820 ;
    END
  END S
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 0.990 1.120 1.650 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.880 1.330 3.080 1.640 ;
        RECT 2.810 0.990 3.080 1.330 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.663100 ;
    PORT
      LAYER li1 ;
        RECT 3.685 1.500 3.855 2.460 ;
        RECT 3.685 1.060 3.960 1.500 ;
        RECT 3.685 0.600 3.855 1.060 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.000 0.345 2.460 ;
        RECT 2.050 2.170 2.680 2.340 ;
        RECT 0.175 1.830 2.070 2.000 ;
        RECT 0.175 1.640 0.345 1.830 ;
        RECT 0.100 1.470 0.345 1.640 ;
        RECT 0.100 0.790 0.270 1.470 ;
        RECT 1.900 0.990 2.070 1.830 ;
        RECT 2.510 1.980 2.680 2.170 ;
        RECT 2.510 1.810 3.510 1.980 ;
        RECT 3.340 0.810 3.510 1.810 ;
        RECT 0.100 0.710 0.350 0.790 ;
        RECT 0.090 0.540 0.350 0.710 ;
        RECT 0.170 0.460 0.350 0.540 ;
        RECT 2.720 0.640 3.510 0.810 ;
        RECT 2.720 0.480 2.890 0.640 ;
        RECT 1.490 0.310 2.890 0.480 ;
  END
END sky130_as_sc_hs__mux2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__mux2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.120 5.520 1.020 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.520 2.810 ;
        RECT 0.650 2.170 0.820 2.630 ;
        RECT 3.095 2.170 3.265 2.630 ;
        RECT 4.115 1.570 4.285 2.630 ;
        RECT 4.975 1.460 5.145 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.280 0.860 0.450 ;
        RECT 3.060 0.300 3.400 0.470 ;
        RECT 0.595 0.105 0.775 0.280 ;
        RECT 3.130 0.105 3.310 0.300 ;
        RECT 4.115 0.105 4.285 0.920 ;
        RECT 4.975 0.105 5.145 0.920 ;
        RECT 0.000 -0.085 5.520 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 1.330 2.560 1.640 ;
        RECT 0.450 0.990 0.720 1.330 ;
        RECT 0.550 0.820 0.720 0.990 ;
        RECT 1.420 0.990 1.620 1.330 ;
        RECT 2.330 0.990 2.570 1.330 ;
        RECT 1.420 0.820 1.590 0.990 ;
        RECT 2.380 0.820 2.550 0.990 ;
        RECT 0.550 0.650 2.550 0.820 ;
    END
  END S
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 0.990 1.120 1.650 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.870 1.330 3.080 1.640 ;
        RECT 2.810 0.990 3.080 1.330 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.122300 ;
    PORT
      LAYER li1 ;
        RECT 3.685 1.500 3.855 2.460 ;
        RECT 3.685 1.380 3.960 1.500 ;
        RECT 4.545 1.380 4.740 2.460 ;
        RECT 3.685 1.210 4.740 1.380 ;
        RECT 3.685 1.060 3.960 1.210 ;
        RECT 3.685 0.600 3.855 1.060 ;
        RECT 4.545 0.600 4.740 1.210 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.000 0.345 2.460 ;
        RECT 2.050 2.170 2.680 2.340 ;
        RECT 0.175 1.830 2.070 2.000 ;
        RECT 0.175 1.640 0.345 1.830 ;
        RECT 0.100 1.470 0.345 1.640 ;
        RECT 0.100 0.790 0.270 1.470 ;
        RECT 1.900 0.990 2.070 1.830 ;
        RECT 2.510 1.980 2.680 2.170 ;
        RECT 2.510 1.810 3.510 1.980 ;
        RECT 3.340 0.810 3.510 1.810 ;
        RECT 0.100 0.710 0.350 0.790 ;
        RECT 0.090 0.540 0.350 0.710 ;
        RECT 0.170 0.460 0.350 0.540 ;
        RECT 2.720 0.640 3.510 0.810 ;
        RECT 2.720 0.480 2.890 0.640 ;
        RECT 1.490 0.310 2.890 0.480 ;
  END
END sky130_as_sc_hs__mux2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 2.300 1.020 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 0.175 1.590 0.345 2.630 ;
        RECT 1.035 1.920 1.205 2.630 ;
        RECT 1.900 1.920 2.070 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.105 0.820 0.540 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.468000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.050 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.468000 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.610 1.340 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.694400 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.750 0.800 2.410 ;
        RECT 1.430 1.750 1.670 2.430 ;
        RECT 0.580 1.530 2.160 1.750 ;
        RECT 1.780 0.890 2.160 1.530 ;
        RECT 1.380 0.710 2.160 0.890 ;
        RECT 1.380 0.620 1.720 0.710 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.150 0.710 1.210 0.880 ;
        RECT 0.150 0.280 0.380 0.710 ;
        RECT 1.000 0.450 1.210 0.710 ;
        RECT 1.870 0.450 2.200 0.540 ;
        RECT 1.000 0.280 2.200 0.450 ;
  END
END sky130_as_sc_hs__nand2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.140 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.175 1.480 0.345 2.630 ;
        RECT 1.035 1.850 1.205 2.630 ;
        RECT 1.895 1.850 2.065 2.630 ;
        RECT 2.755 1.850 2.925 2.630 ;
        RECT 3.615 1.470 3.785 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.530 ;
        RECT 1.465 0.105 1.635 0.530 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.400 1.040 1.840 1.310 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 2.120 1.040 3.010 1.310 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.472800 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.680 0.775 2.460 ;
        RECT 1.465 1.680 1.635 2.460 ;
        RECT 2.325 1.680 2.495 2.460 ;
        RECT 3.185 1.680 3.355 2.460 ;
        RECT 0.605 1.510 3.435 1.680 ;
        RECT 3.185 0.860 3.435 1.510 ;
        RECT 2.235 0.690 3.440 0.860 ;
        RECT 2.235 0.680 2.575 0.690 ;
        RECT 3.100 0.670 3.440 0.690 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 0.700 2.065 0.870 ;
        RECT 0.175 0.280 0.345 0.700 ;
        RECT 1.035 0.280 1.205 0.700 ;
        RECT 1.895 0.450 2.065 0.700 ;
        RECT 3.615 0.450 3.785 0.930 ;
        RECT 1.895 0.280 3.785 0.450 ;
  END
END sky130_as_sc_hs__nand2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 3.680 1.020 ;
        RECT 0.130 -0.075 0.380 0.110 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
        RECT 1.510 -0.100 1.830 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.300 0.105 0.540 0.830 ;
        RECT 1.940 0.105 2.200 0.540 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.300 1.650 0.540 2.630 ;
        RECT 1.280 1.600 1.520 2.630 ;
        RECT 2.190 1.920 2.600 2.630 ;
        RECT 3.250 1.920 3.480 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    PORT
      LAYER li1 ;
        RECT 3.280 1.370 3.460 1.750 ;
        RECT 3.150 1.040 3.460 1.370 ;
        RECT 3.280 0.840 3.460 1.040 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699800 ;
    PORT
      LAYER li1 ;
        RECT 1.720 1.750 1.960 2.430 ;
        RECT 2.810 1.750 3.050 2.430 ;
        RECT 1.720 1.530 3.050 1.750 ;
        RECT 2.370 1.270 2.610 1.530 ;
        RECT 2.370 1.050 2.980 1.270 ;
        RECT 2.760 0.870 2.980 1.050 ;
        RECT 2.760 0.620 3.100 0.870 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.250 1.060 0.600 1.400 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.770 1.340 1.000 2.460 ;
        RECT 0.770 1.050 2.200 1.340 ;
        RECT 0.770 0.290 1.000 1.050 ;
        RECT 1.530 0.710 2.590 0.880 ;
        RECT 1.530 0.280 1.760 0.710 ;
        RECT 2.380 0.450 2.590 0.710 ;
        RECT 3.250 0.450 3.580 0.540 ;
        RECT 2.380 0.280 3.580 0.450 ;
  END
END sky130_as_sc_hs__nand2b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand3_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.100 3.680 1.020 ;
        RECT 0.130 -0.100 0.450 0.100 ;
        RECT 2.430 -0.075 2.680 0.100 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.175 1.590 0.345 2.630 ;
        RECT 1.035 1.920 1.205 2.630 ;
        RECT 1.900 2.180 2.610 2.630 ;
        RECT 3.325 1.920 3.495 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.105 0.820 0.540 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.050 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.610 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.489000 ;
    PORT
      LAYER li1 ;
        RECT 2.280 1.340 2.470 1.670 ;
        RECT 2.210 1.080 2.630 1.340 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008000 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.750 0.800 2.410 ;
        RECT 1.430 2.010 1.670 2.430 ;
        RECT 2.860 2.010 3.100 2.430 ;
        RECT 1.430 1.840 3.100 2.010 ;
        RECT 1.430 1.750 1.670 1.840 ;
        RECT 0.580 1.530 1.670 1.750 ;
        RECT 2.860 0.890 3.100 1.840 ;
        RECT 2.810 0.620 3.150 0.890 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.150 0.710 1.210 0.880 ;
        RECT 0.150 0.280 0.380 0.710 ;
        RECT 1.000 0.450 1.210 0.710 ;
        RECT 1.380 0.680 2.630 0.890 ;
        RECT 1.380 0.620 1.720 0.680 ;
        RECT 1.850 0.450 2.180 0.510 ;
        RECT 1.000 0.280 2.180 0.450 ;
        RECT 2.420 0.450 2.630 0.680 ;
        RECT 3.315 0.450 3.580 0.570 ;
        RECT 2.420 0.280 3.580 0.450 ;
  END
END sky130_as_sc_hs__nand3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand4_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 4.600 1.020 ;
        RECT 0.000 0.100 3.680 0.130 ;
        RECT 0.130 -0.100 0.450 0.100 ;
        RECT 2.430 -0.075 2.680 0.100 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.175 1.590 0.345 2.630 ;
        RECT 1.035 1.920 1.205 2.630 ;
        RECT 1.900 2.180 2.610 2.630 ;
        RECT 3.310 2.170 3.510 2.630 ;
        RECT 4.185 1.930 4.355 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.105 0.820 0.540 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.489000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.050 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.489000 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.810 1.290 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.489000 ;
    PORT
      LAYER li1 ;
        RECT 2.280 1.280 2.480 1.670 ;
        RECT 2.210 1.060 2.630 1.280 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.283800 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.750 0.800 2.410 ;
        RECT 1.430 2.010 1.670 2.430 ;
        RECT 2.860 2.010 3.100 2.110 ;
        RECT 1.430 2.000 3.100 2.010 ;
        RECT 3.740 2.000 3.940 2.280 ;
        RECT 1.430 1.840 3.940 2.000 ;
        RECT 1.430 1.750 1.670 1.840 ;
        RECT 2.860 1.830 3.940 1.840 ;
        RECT 0.580 1.580 1.670 1.750 ;
        RECT 3.740 1.760 3.940 1.830 ;
        RECT 3.740 1.580 4.230 1.760 ;
        RECT 3.980 0.880 4.230 1.580 ;
        RECT 3.675 0.680 4.230 0.880 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.489000 ;
    PORT
      LAYER li1 ;
        RECT 3.360 1.340 3.560 1.660 ;
        RECT 3.360 1.060 3.810 1.340 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.150 0.710 1.210 0.880 ;
        RECT 0.150 0.280 0.380 0.710 ;
        RECT 1.000 0.450 1.210 0.710 ;
        RECT 1.380 0.670 3.145 0.890 ;
        RECT 1.850 0.450 2.180 0.480 ;
        RECT 1.000 0.280 2.180 0.450 ;
        RECT 2.350 0.450 2.710 0.480 ;
        RECT 3.315 0.450 3.505 0.620 ;
        RECT 4.050 0.450 4.435 0.510 ;
        RECT 2.350 0.280 4.435 0.450 ;
  END
END sky130_as_sc_hs__nand4_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.020 2.300 1.020 ;
        RECT 0.130 -0.100 0.450 -0.020 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 0.550 1.970 0.830 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.860 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.900 0.105 2.070 0.540 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.390 1.060 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.610 1.340 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641200 ;
    PORT
      LAYER li1 ;
        RECT 1.460 1.750 1.640 1.860 ;
        RECT 1.460 1.520 2.160 1.750 ;
        RECT 1.870 0.890 2.160 1.520 ;
        RECT 0.600 0.710 2.160 0.890 ;
        RECT 0.600 0.520 0.780 0.710 ;
        RECT 1.460 0.500 1.640 0.710 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.170 1.740 0.350 2.460 ;
        RECT 1.030 2.290 2.100 2.460 ;
        RECT 1.030 1.740 1.210 2.290 ;
        RECT 1.930 2.130 2.100 2.290 ;
        RECT 0.170 1.570 1.210 1.740 ;
  END
END sky130_as_sc_hs__nor2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.140 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.605 1.850 0.775 2.630 ;
        RECT 1.465 1.850 1.635 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.870 ;
        RECT 0.950 0.290 1.290 0.510 ;
        RECT 1.810 0.290 2.150 0.510 ;
        RECT 2.670 0.290 3.010 0.510 ;
        RECT 1.035 0.105 1.205 0.290 ;
        RECT 1.895 0.105 2.065 0.290 ;
        RECT 2.755 0.105 2.925 0.290 ;
        RECT 3.625 0.105 3.795 0.930 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 0.400 1.040 1.840 1.310 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.984000 ;
    PORT
      LAYER li1 ;
        RECT 2.120 1.040 3.010 1.310 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.282400 ;
    PORT
      LAYER li1 ;
        RECT 2.240 1.740 2.560 1.770 ;
        RECT 3.130 1.740 3.435 1.820 ;
        RECT 2.240 1.570 3.435 1.740 ;
        RECT 2.240 1.550 2.560 1.570 ;
        RECT 3.130 1.500 3.435 1.570 ;
        RECT 3.185 0.850 3.435 1.500 ;
        RECT 0.520 0.680 3.435 0.850 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.680 0.345 2.450 ;
        RECT 1.035 1.680 1.205 2.450 ;
        RECT 1.895 2.280 3.795 2.450 ;
        RECT 1.895 1.680 2.065 2.280 ;
        RECT 2.755 2.000 2.925 2.280 ;
        RECT 0.175 1.510 2.065 1.680 ;
        RECT 3.625 1.450 3.795 2.280 ;
  END
END sky130_as_sc_hs__nor2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.100 3.680 1.020 ;
        RECT 0.130 -0.100 0.450 0.100 ;
        RECT 2.430 -0.075 2.680 0.100 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.550 1.970 0.830 2.630 ;
        RECT 3.270 1.590 3.460 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.860 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.900 0.105 2.070 0.830 ;
        RECT 3.280 0.105 3.450 0.830 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.060 0.980 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641200 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.400 1.680 2.070 ;
        RECT 1.150 1.210 1.680 1.400 ;
        RECT 1.150 0.890 1.380 1.210 ;
        RECT 0.570 0.710 1.660 0.890 ;
        RECT 0.570 0.280 0.790 0.710 ;
        RECT 1.440 0.280 1.660 0.710 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.230 1.000 3.530 1.420 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 0.150 1.800 0.380 2.460 ;
        RECT 1.000 2.240 2.130 2.460 ;
        RECT 1.000 1.800 1.240 2.240 ;
        RECT 1.850 1.920 2.130 2.240 ;
        RECT 0.150 1.570 1.240 1.800 ;
        RECT 1.870 1.240 2.080 1.360 ;
        RECT 2.810 1.240 3.060 2.430 ;
        RECT 1.870 1.020 3.060 1.240 ;
        RECT 1.870 1.000 2.080 1.020 ;
        RECT 2.810 0.280 3.060 1.020 ;
  END
END sky130_as_sc_hs__nor2b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor3_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.100 3.680 1.020 ;
        RECT 0.130 -0.100 0.450 0.100 ;
        RECT 2.430 -0.075 2.680 0.100 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.570 2.060 0.810 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.920 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.900 0.105 2.650 0.540 ;
        RECT 3.325 0.105 3.495 0.910 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.490500 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.090 0.930 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.490500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 1.060 1.870 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.490500 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.310 2.280 1.610 ;
        RECT 2.110 1.090 2.630 1.310 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.821800 ;
    PORT
      LAYER li1 ;
        RECT 2.870 1.460 3.080 1.790 ;
        RECT 2.870 0.880 3.100 1.460 ;
        RECT 0.605 0.870 3.100 0.880 ;
        RECT 0.605 0.710 3.065 0.870 ;
        RECT 0.605 0.460 0.775 0.710 ;
        RECT 1.465 0.410 1.635 0.710 ;
        RECT 2.895 0.510 3.065 0.710 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.160 1.890 0.360 2.450 ;
        RECT 1.020 2.280 2.080 2.450 ;
        RECT 1.020 1.890 1.215 2.280 ;
        RECT 1.880 2.120 2.080 2.280 ;
        RECT 2.450 2.020 3.520 2.210 ;
        RECT 2.450 1.950 2.650 2.020 ;
        RECT 0.160 1.720 1.215 1.890 ;
        RECT 1.385 1.780 2.650 1.950 ;
        RECT 2.450 1.510 2.650 1.780 ;
        RECT 3.320 1.490 3.520 2.020 ;
  END
END sky130_as_sc_hs__nor3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oa21_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oa21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 3.680 1.020 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 1.035 2.190 1.205 2.630 ;
        RECT 2.225 1.550 2.395 2.630 ;
        RECT 3.085 1.550 3.255 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.280 0.860 0.450 ;
        RECT 0.605 0.105 0.775 0.280 ;
        RECT 2.225 0.105 2.395 0.820 ;
        RECT 3.085 0.105 3.255 0.900 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.260 0.990 0.550 1.380 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.810 0.990 1.050 1.680 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 0.990 1.510 1.670 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 2.655 1.490 2.825 2.460 ;
        RECT 2.650 0.950 2.900 1.490 ;
        RECT 2.655 0.480 2.825 0.950 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.020 0.345 2.290 ;
        RECT 1.680 2.020 1.850 2.460 ;
        RECT 0.175 1.850 1.850 2.020 ;
        RECT 0.175 1.550 0.345 1.850 ;
        RECT 1.680 1.250 1.850 1.850 ;
        RECT 2.180 1.250 2.350 1.330 ;
        RECT 1.680 1.080 2.350 1.250 ;
        RECT 0.175 0.650 1.205 0.820 ;
        RECT 0.175 0.450 0.345 0.650 ;
        RECT 1.035 0.430 1.205 0.650 ;
        RECT 1.680 0.550 1.850 1.080 ;
        RECT 2.180 1.000 2.350 1.080 ;
  END
END sky130_as_sc_hs__oa21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oa21_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oa21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.150 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 1.035 2.190 1.205 2.630 ;
        RECT 2.225 1.550 2.395 2.630 ;
        RECT 3.085 1.550 3.255 2.630 ;
        RECT 3.945 1.550 4.115 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.280 0.860 0.450 ;
        RECT 0.605 0.105 0.775 0.280 ;
        RECT 2.225 0.105 2.395 0.820 ;
        RECT 3.085 0.105 3.255 0.900 ;
        RECT 3.945 0.105 4.115 0.900 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.260 0.990 0.550 1.380 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.810 0.990 1.050 1.680 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 0.990 1.510 1.670 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 2.655 1.490 2.825 2.460 ;
        RECT 2.650 1.330 2.880 1.490 ;
        RECT 3.515 1.330 3.685 2.460 ;
        RECT 2.650 1.090 3.685 1.330 ;
        RECT 2.650 0.950 2.880 1.090 ;
        RECT 2.655 0.600 2.825 0.950 ;
        RECT 3.515 0.490 3.685 1.090 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.020 0.345 2.240 ;
        RECT 1.680 2.020 1.850 2.460 ;
        RECT 0.175 1.850 1.850 2.020 ;
        RECT 0.175 1.550 0.345 1.850 ;
        RECT 1.680 1.250 1.850 1.850 ;
        RECT 2.180 1.250 2.350 1.330 ;
        RECT 1.680 1.080 2.350 1.250 ;
        RECT 0.175 0.650 1.205 0.820 ;
        RECT 0.175 0.490 0.345 0.650 ;
        RECT 1.035 0.490 1.205 0.650 ;
        RECT 1.680 0.520 1.850 1.080 ;
        RECT 2.180 1.000 2.350 1.080 ;
  END
END sky130_as_sc_hs__oa21_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oa22_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oa22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.140 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.175 2.140 0.345 2.630 ;
        RECT 2.230 1.590 2.960 2.630 ;
        RECT 3.645 1.610 3.815 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.290 0.860 0.460 ;
        RECT 2.700 0.290 3.040 0.460 ;
        RECT 0.605 0.105 0.775 0.290 ;
        RECT 2.785 0.105 2.955 0.290 ;
        RECT 3.645 0.105 3.815 0.830 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 1.330 0.440 1.970 ;
        RECT 0.190 1.000 0.550 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.330 0.930 1.910 ;
        RECT 0.720 1.000 1.030 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 1.330 1.450 1.880 ;
        RECT 1.200 1.000 1.510 1.330 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.020 0.970 2.450 1.420 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 3.215 1.470 3.385 2.460 ;
        RECT 3.215 0.970 3.540 1.470 ;
        RECT 3.215 0.280 3.385 0.970 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.035 2.220 1.205 2.460 ;
        RECT 1.035 2.050 1.850 2.220 ;
        RECT 1.680 0.830 1.850 2.050 ;
        RECT 0.175 0.660 1.205 0.830 ;
        RECT 0.175 0.280 0.345 0.660 ;
        RECT 1.035 0.450 1.205 0.660 ;
        RECT 1.430 0.800 1.850 0.830 ;
        RECT 2.720 1.000 3.040 1.340 ;
        RECT 2.720 0.800 2.890 1.000 ;
        RECT 1.430 0.630 2.890 0.800 ;
        RECT 1.035 0.280 2.475 0.450 ;
  END
END sky130_as_sc_hs__oa22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oa22_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oa22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 5.060 1.020 ;
        RECT 0.000 0.140 4.140 0.150 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.060 2.810 ;
        RECT 0.175 2.140 0.345 2.630 ;
        RECT 2.230 1.590 2.960 2.630 ;
        RECT 3.645 1.610 3.815 2.630 ;
        RECT 4.505 1.460 4.675 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.290 0.860 0.460 ;
        RECT 2.700 0.290 3.040 0.460 ;
        RECT 0.605 0.105 0.775 0.290 ;
        RECT 2.785 0.105 2.955 0.290 ;
        RECT 3.645 0.105 3.815 0.830 ;
        RECT 4.505 0.105 4.675 0.960 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 1.330 0.440 1.970 ;
        RECT 0.190 1.000 0.550 1.330 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.330 0.930 1.910 ;
        RECT 0.720 1.000 1.030 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 1.330 1.450 1.880 ;
        RECT 1.200 1.000 1.510 1.330 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.020 0.970 2.450 1.420 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 3.215 1.470 3.385 2.460 ;
        RECT 3.215 1.350 3.540 1.470 ;
        RECT 4.075 1.350 4.245 2.460 ;
        RECT 3.215 1.050 4.245 1.350 ;
        RECT 3.215 0.970 3.540 1.050 ;
        RECT 3.215 0.280 3.385 0.970 ;
        RECT 4.075 0.280 4.245 1.050 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 1.035 2.220 1.205 2.460 ;
        RECT 1.035 2.050 1.850 2.220 ;
        RECT 1.680 0.830 1.850 2.050 ;
        RECT 0.175 0.660 1.205 0.830 ;
        RECT 0.175 0.280 0.345 0.660 ;
        RECT 1.035 0.450 1.205 0.660 ;
        RECT 1.430 0.800 1.850 0.830 ;
        RECT 2.720 1.000 3.040 1.340 ;
        RECT 2.720 0.800 2.890 1.000 ;
        RECT 1.430 0.630 2.890 0.800 ;
        RECT 1.035 0.280 2.475 0.450 ;
  END
END sky130_as_sc_hs__oa22_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oai21_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oai21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 3.220 1.020 ;
        RECT 0.000 0.110 2.300 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.220 2.810 ;
        RECT 0.175 1.880 0.345 2.630 ;
        RECT 1.895 2.180 2.065 2.630 ;
        RECT 2.755 2.180 2.925 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.280 0.860 0.450 ;
        RECT 1.380 0.280 1.720 0.450 ;
        RECT 0.605 0.105 0.775 0.280 ;
        RECT 1.465 0.105 1.635 0.280 ;
        RECT 0.000 -0.085 3.220 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.220 1.500 1.860 1.670 ;
        RECT 0.220 0.990 0.470 1.500 ;
        RECT 1.620 1.350 1.860 1.500 ;
        RECT 1.620 0.990 1.890 1.350 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.830 1.010 1.410 1.330 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.100 1.350 2.330 1.670 ;
        RECT 2.100 0.990 2.370 1.350 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.736400 ;
    PORT
      LAYER li1 ;
        RECT 2.325 2.010 2.495 2.460 ;
        RECT 0.955 1.840 2.710 2.010 ;
        RECT 2.540 1.740 2.710 1.840 ;
        RECT 2.540 1.000 2.830 1.740 ;
        RECT 2.540 0.810 2.710 1.000 ;
        RECT 2.240 0.640 2.710 0.810 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.520 2.270 1.725 2.440 ;
        RECT 0.175 0.650 2.065 0.820 ;
        RECT 0.175 0.280 0.345 0.650 ;
        RECT 1.035 0.280 1.205 0.650 ;
        RECT 1.895 0.450 2.065 0.650 ;
        RECT 1.895 0.280 3.010 0.450 ;
  END
END sky130_as_sc_hs__oai21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__oai22_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__oai22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.140 4.600 1.020 ;
        RECT 0.000 0.110 3.680 0.140 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.600 2.810 ;
        RECT 0.615 2.140 0.785 2.630 ;
        RECT 3.735 1.940 3.905 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.770 0.300 3.120 0.490 ;
        RECT 3.640 0.300 3.995 0.490 ;
        RECT 2.865 0.105 3.035 0.300 ;
        RECT 3.735 0.105 3.905 0.300 ;
        RECT 0.000 -0.085 4.600 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.360 0.650 1.530 ;
        RECT 0.310 1.020 0.990 1.360 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 1.160 1.020 1.620 1.360 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 2.650 1.020 3.220 1.360 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 3.530 1.020 4.020 1.360 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928300 ;
    PORT
      LAYER li1 ;
        RECT 1.475 1.770 1.645 2.120 ;
        RECT 2.865 1.770 3.035 2.120 ;
        RECT 1.390 1.600 3.120 1.770 ;
        RECT 1.790 0.840 2.160 1.600 ;
        RECT 0.520 0.670 2.160 0.840 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.180 1.870 0.360 2.460 ;
        RECT 1.045 2.290 2.075 2.460 ;
        RECT 1.045 1.870 1.215 2.290 ;
        RECT 1.905 1.940 2.075 2.290 ;
        RECT 2.425 2.290 3.475 2.460 ;
        RECT 2.425 1.940 2.595 2.290 ;
        RECT 0.180 1.700 1.215 1.870 ;
        RECT 3.305 1.770 3.475 2.290 ;
        RECT 4.165 1.770 4.335 2.460 ;
        RECT 3.305 1.600 4.335 1.770 ;
        RECT 0.175 0.450 0.345 0.840 ;
        RECT 4.165 0.830 4.335 0.900 ;
        RECT 2.410 0.660 4.335 0.830 ;
        RECT 2.410 0.450 2.580 0.660 ;
        RECT 0.175 0.280 2.580 0.450 ;
        RECT 3.295 0.280 3.465 0.660 ;
        RECT 4.165 0.290 4.335 0.660 ;
  END
END sky130_as_sc_hs__oai22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__or2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 2.300 1.020 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 1.035 1.950 1.205 2.630 ;
        RECT 1.875 2.250 2.210 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 0.955 0.305 1.285 0.475 ;
        RECT 1.035 0.105 1.205 0.305 ;
        RECT 1.875 0.300 2.210 0.490 ;
        RECT 1.955 0.105 2.125 0.300 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.390 1.430 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.760 0.990 1.010 1.440 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.459200 ;
    PORT
      LAYER li1 ;
        RECT 1.525 2.080 1.695 2.280 ;
        RECT 1.525 1.950 1.970 2.080 ;
        RECT 1.560 1.910 1.970 1.950 ;
        RECT 1.720 0.860 1.970 1.910 ;
        RECT 1.700 0.830 1.970 0.860 ;
        RECT 1.525 0.770 1.970 0.830 ;
        RECT 1.525 0.660 1.870 0.770 ;
        RECT 1.525 0.420 1.695 0.660 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.780 0.345 2.460 ;
        RECT 0.175 1.610 1.450 1.780 ;
        RECT 0.175 1.600 0.530 1.610 ;
        RECT 1.280 1.400 1.450 1.610 ;
        RECT 1.185 1.330 1.450 1.400 ;
        RECT 1.185 1.000 1.550 1.330 ;
        RECT 1.185 0.820 1.355 1.000 ;
        RECT 0.560 0.650 1.355 0.820 ;
        RECT 0.560 0.450 0.775 0.650 ;
  END
END sky130_as_sc_hs__or2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__or2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 3.220 1.020 ;
        RECT 0.000 0.110 2.300 0.130 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.220 2.810 ;
        RECT 1.035 1.950 1.205 2.630 ;
        RECT 1.890 2.250 2.230 2.630 ;
        RECT 2.835 1.430 3.005 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.830 ;
        RECT 1.035 0.105 1.205 0.830 ;
        RECT 1.890 0.300 2.230 0.490 ;
        RECT 1.955 0.105 2.125 0.300 ;
        RECT 2.835 0.105 3.005 0.910 ;
        RECT 0.000 -0.085 3.220 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.170 1.000 0.400 1.430 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 1.000 1.130 1.440 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.918400 ;
    PORT
      LAYER li1 ;
        RECT 1.515 2.080 1.715 2.280 ;
        RECT 1.515 1.950 1.960 2.080 ;
        RECT 1.570 1.910 1.960 1.950 ;
        RECT 1.730 1.270 1.960 1.910 ;
        RECT 2.405 1.270 2.580 2.460 ;
        RECT 1.730 1.100 2.580 1.270 ;
        RECT 1.730 0.830 1.940 1.100 ;
        RECT 1.515 0.770 1.940 0.830 ;
        RECT 1.515 0.660 1.900 0.770 ;
        RECT 1.515 0.450 1.715 0.660 ;
        RECT 2.400 0.600 2.580 1.100 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.780 0.345 2.460 ;
        RECT 0.175 1.740 1.460 1.780 ;
        RECT 0.175 1.610 1.475 1.740 ;
        RECT 0.175 1.600 0.740 1.610 ;
        RECT 0.570 0.860 0.740 1.600 ;
        RECT 1.305 1.330 1.475 1.610 ;
        RECT 1.305 1.000 1.560 1.330 ;
        RECT 0.570 0.450 0.775 0.860 ;
  END
END sky130_as_sc_hs__or2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__pulsed_dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__pulsed_dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.170 11.960 1.020 ;
        RECT 0.000 0.160 8.280 0.170 ;
        RECT 10.110 0.160 11.500 0.170 ;
        RECT 0.000 0.120 7.360 0.160 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 5.495 0.110 5.520 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 11.960 2.810 ;
        RECT 0.810 1.570 0.980 2.630 ;
        RECT 2.415 1.580 2.585 2.630 ;
        RECT 4.485 2.040 4.655 2.630 ;
        RECT 5.775 1.510 5.945 2.630 ;
        RECT 8.695 2.180 8.865 2.630 ;
        RECT 10.265 1.510 10.435 2.630 ;
        RECT 11.280 1.450 11.450 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.760 0.280 1.090 0.450 ;
        RECT 2.330 0.280 2.670 0.450 ;
        RECT 3.450 0.300 3.790 0.470 ;
        RECT 4.400 0.300 4.740 0.470 ;
        RECT 5.690 0.300 6.030 0.470 ;
        RECT 8.610 0.300 8.950 0.470 ;
        RECT 0.840 0.105 1.010 0.280 ;
        RECT 2.415 0.105 2.585 0.280 ;
        RECT 3.535 0.105 3.705 0.300 ;
        RECT 4.485 0.105 4.655 0.300 ;
        RECT 5.775 0.105 5.945 0.300 ;
        RECT 8.695 0.105 8.865 0.300 ;
        RECT 10.265 0.105 10.435 0.540 ;
        RECT 11.280 0.105 11.450 0.930 ;
        RECT 0.000 -0.085 11.960 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.520 0.980 0.790 1.330 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 5.660 0.980 5.930 1.330 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.688800 ;
    PORT
      LAYER li1 ;
        RECT 10.820 1.540 10.990 2.460 ;
        RECT 10.820 0.820 11.090 1.540 ;
        RECT 10.820 0.570 10.990 0.820 ;
    END
  END Q
  PIN PULSE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.507800 ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.700 3.705 2.460 ;
        RECT 3.535 1.530 4.960 1.700 ;
        RECT 3.965 0.600 4.135 1.530 ;
        RECT 4.790 0.980 4.960 1.530 ;
        RECT 6.550 0.980 6.720 1.330 ;
        RECT 8.010 0.980 8.180 1.330 ;
      LAYER met1 ;
        RECT 6.450 2.210 8.180 2.220 ;
        RECT 4.310 2.040 8.180 2.210 ;
        RECT 4.310 1.730 4.480 2.040 ;
        RECT 4.280 1.470 4.510 1.730 ;
        RECT 6.550 1.290 6.720 2.040 ;
        RECT 8.010 1.330 8.180 2.040 ;
        RECT 6.520 1.020 6.750 1.290 ;
        RECT 7.970 1.020 8.220 1.330 ;
    END
  END PULSE
  PIN PULSEN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    ANTENNADIFFAREA 0.738000 ;
    PORT
      LAYER li1 ;
        RECT 5.130 0.580 5.300 2.460 ;
        RECT 7.030 0.980 7.200 1.330 ;
      LAYER met1 ;
        RECT 7.000 1.050 7.230 1.320 ;
        RECT 5.100 0.600 5.330 0.890 ;
        RECT 7.030 0.600 7.200 1.050 ;
        RECT 5.100 0.430 7.200 0.600 ;
    END
  END PULSEN
  OBS
      LAYER li1 ;
        RECT 0.175 0.810 0.345 2.460 ;
        RECT 1.440 1.330 1.610 2.460 ;
        RECT 1.050 0.810 1.220 1.330 ;
        RECT 0.175 0.640 1.220 0.810 ;
        RECT 1.440 0.980 1.810 1.330 ;
        RECT 1.985 1.250 2.155 2.460 ;
        RECT 2.960 1.340 3.130 2.460 ;
        RECT 2.620 1.250 2.790 1.340 ;
        RECT 1.985 1.080 2.790 1.250 ;
        RECT 0.175 0.580 0.345 0.640 ;
        RECT 1.440 0.580 1.610 0.980 ;
        RECT 1.985 0.580 2.155 1.080 ;
        RECT 2.620 0.990 2.790 1.080 ;
        RECT 2.960 0.990 3.390 1.340 ;
        RECT 2.960 0.580 3.130 0.990 ;
        RECT 4.310 0.980 4.480 1.330 ;
        RECT 6.205 0.570 6.375 2.460 ;
        RECT 7.370 0.810 7.540 2.460 ;
        RECT 9.310 1.770 9.480 2.460 ;
        RECT 8.490 1.600 9.480 1.770 ;
        RECT 8.490 0.980 8.660 1.600 ;
        RECT 9.310 1.340 9.480 1.600 ;
        RECT 8.970 0.810 9.140 1.330 ;
        RECT 7.370 0.640 9.140 0.810 ;
        RECT 9.310 0.990 9.620 1.340 ;
        RECT 9.835 1.250 10.005 2.460 ;
        RECT 10.420 1.250 10.650 1.340 ;
        RECT 9.835 1.080 10.650 1.250 ;
        RECT 7.370 0.570 7.540 0.640 ;
        RECT 9.310 0.570 9.480 0.990 ;
        RECT 9.835 0.570 10.005 1.080 ;
        RECT 10.420 0.990 10.650 1.080 ;
      LAYER met1 ;
        RECT 4.280 0.980 4.510 1.310 ;
        RECT 0.990 0.810 1.380 0.840 ;
        RECT 4.310 0.810 4.480 0.980 ;
        RECT 0.990 0.640 4.480 0.810 ;
        RECT 0.990 0.610 1.380 0.640 ;
  END
END sky130_as_sc_hs__pulsed_dfxtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tap_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
        RECT 0.110 1.460 0.340 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.110 0.460 1.020 ;
        RECT 0.090 -0.120 0.400 0.110 ;
      LAYER li1 ;
        RECT 0.120 0.105 0.340 1.000 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__tap_1


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tieh
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.730 1.840 1.040 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 0.380 1.040 1.630 ;
    END
  END ONE
END sky130_as_sc_hs__tieh


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tiel
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.105 1.040 0.860 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ZERO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 1.140 1.040 2.390 ;
    END
  END ZERO
END sky130_as_sc_hs__tiel


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 5.060 1.020 ;
        RECT 0.000 0.120 4.600 0.130 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 3.910 0.110 4.060 0.120 ;
        RECT 4.435 0.110 4.585 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.060 2.810 ;
        RECT 0.605 2.060 0.775 2.630 ;
        RECT 3.580 2.190 3.750 2.630 ;
        RECT 4.690 1.610 4.860 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.590 ;
        RECT 3.590 0.105 3.760 0.830 ;
        RECT 4.640 0.105 4.810 0.540 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.409500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.680 1.220 1.850 ;
        RECT 0.445 1.100 0.680 1.680 ;
        RECT 2.720 1.000 2.940 1.330 ;
        RECT 2.720 0.900 2.890 1.000 ;
        RECT 2.130 0.730 2.890 0.900 ;
        RECT 2.130 0.660 2.300 0.730 ;
      LAYER met1 ;
        RECT 0.990 1.640 1.410 1.910 ;
        RECT 1.240 0.910 1.410 1.640 ;
        RECT 1.240 0.730 2.360 0.910 ;
        RECT 2.070 0.630 2.360 0.730 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615000 ;
    PORT
      LAYER li1 ;
        RECT 4.210 1.780 4.380 2.430 ;
        RECT 4.210 1.530 4.470 1.780 ;
        RECT 4.300 1.500 4.470 1.530 ;
        RECT 4.300 0.900 4.560 1.500 ;
        RECT 4.300 0.830 4.470 0.900 ;
        RECT 4.210 0.650 4.470 0.830 ;
        RECT 4.210 0.500 4.380 0.650 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.460 1.000 3.700 1.330 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 0.100 2.020 0.345 2.440 ;
        RECT 1.390 2.060 3.410 2.230 ;
        RECT 0.100 0.930 0.275 2.020 ;
        RECT 0.880 1.040 1.210 1.260 ;
        RECT 0.880 0.930 1.050 1.040 ;
        RECT 0.100 0.760 1.050 0.930 ;
        RECT 1.390 0.830 1.560 2.060 ;
        RECT 3.240 2.010 3.410 2.060 ;
        RECT 3.240 1.840 4.040 2.010 ;
        RECT 2.360 1.670 3.080 1.730 ;
        RECT 1.790 1.500 3.290 1.670 ;
        RECT 1.790 1.330 1.960 1.500 ;
        RECT 1.730 1.000 1.960 1.330 ;
        RECT 2.170 1.070 2.510 1.300 ;
        RECT 0.100 0.750 0.345 0.760 ;
        RECT 0.175 0.280 0.345 0.750 ;
        RECT 1.390 0.640 1.815 0.830 ;
        RECT 1.645 0.450 1.815 0.640 ;
        RECT 3.120 0.560 3.290 1.500 ;
        RECT 3.870 1.330 4.040 1.840 ;
        RECT 3.870 1.000 4.130 1.330 ;
        RECT 1.645 0.280 2.190 0.450 ;
      LAYER met1 ;
        RECT 0.110 2.270 0.400 2.290 ;
        RECT 0.110 2.080 2.330 2.270 ;
        RECT 0.110 2.060 0.400 2.080 ;
        RECT 2.170 1.280 2.330 2.080 ;
        RECT 2.110 1.050 2.400 1.280 ;
  END
END sky130_as_sc_hs__xnor2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.130 5.980 1.020 ;
        RECT 0.000 0.120 4.600 0.130 ;
        RECT 4.650 0.120 5.980 0.130 ;
        RECT 0.000 0.110 3.680 0.120 ;
        RECT 3.910 0.110 4.060 0.120 ;
        RECT 4.520 0.110 4.670 0.120 ;
        RECT 4.950 0.110 5.100 0.120 ;
        RECT 5.380 0.110 5.530 0.120 ;
        RECT 0.130 -0.100 0.450 0.110 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.980 2.810 ;
        RECT 0.605 2.060 0.775 2.630 ;
        RECT 3.580 2.190 3.750 2.630 ;
        RECT 4.725 1.520 4.895 2.630 ;
        RECT 5.585 1.480 5.755 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.590 ;
        RECT 3.590 0.105 3.760 0.830 ;
        RECT 4.725 0.105 4.895 0.900 ;
        RECT 5.585 0.105 5.755 0.900 ;
        RECT 0.000 -0.085 5.980 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.409500 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.680 1.220 1.850 ;
        RECT 0.445 1.100 0.680 1.680 ;
        RECT 2.720 1.000 2.950 1.330 ;
        RECT 2.720 0.900 2.890 1.000 ;
        RECT 2.130 0.730 2.890 0.900 ;
        RECT 2.130 0.660 2.300 0.730 ;
      LAYER met1 ;
        RECT 0.990 1.640 1.410 1.910 ;
        RECT 1.240 0.910 1.410 1.640 ;
        RECT 1.240 0.730 2.360 0.910 ;
        RECT 2.070 0.630 2.360 0.730 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.213600 ;
    PORT
      LAYER li1 ;
        RECT 4.290 1.530 4.470 2.430 ;
        RECT 4.300 1.340 4.540 1.530 ;
        RECT 5.155 1.340 5.325 2.450 ;
        RECT 4.300 1.130 5.325 1.340 ;
        RECT 4.300 0.910 4.540 1.130 ;
        RECT 4.290 0.580 4.470 0.910 ;
        RECT 5.155 0.600 5.325 1.130 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.460 1.000 3.700 1.330 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 0.100 2.020 0.345 2.440 ;
        RECT 1.390 2.060 3.410 2.230 ;
        RECT 0.100 0.930 0.275 2.020 ;
        RECT 0.880 1.040 1.210 1.260 ;
        RECT 0.880 0.930 1.050 1.040 ;
        RECT 0.100 0.760 1.050 0.930 ;
        RECT 1.390 0.830 1.560 2.060 ;
        RECT 3.240 2.010 3.410 2.060 ;
        RECT 3.240 1.840 4.040 2.010 ;
        RECT 2.360 1.670 3.080 1.730 ;
        RECT 1.790 1.500 3.290 1.670 ;
        RECT 1.790 1.330 1.960 1.500 ;
        RECT 1.730 1.000 1.960 1.330 ;
        RECT 2.170 1.070 2.510 1.300 ;
        RECT 0.100 0.750 0.345 0.760 ;
        RECT 0.175 0.280 0.345 0.750 ;
        RECT 1.390 0.640 1.815 0.830 ;
        RECT 1.645 0.450 1.815 0.640 ;
        RECT 3.120 0.490 3.290 1.500 ;
        RECT 3.870 1.330 4.040 1.840 ;
        RECT 3.870 1.000 4.130 1.330 ;
        RECT 1.645 0.280 2.180 0.450 ;
      LAYER met1 ;
        RECT 0.110 2.270 0.400 2.290 ;
        RECT 0.110 2.080 2.330 2.270 ;
        RECT 0.110 2.060 0.400 2.080 ;
        RECT 2.170 1.280 2.330 2.080 ;
        RECT 2.110 1.050 2.400 1.280 ;
  END
END sky130_as_sc_hs__xnor2_4


END LIBRARY
