magic
tech sky130A
magscale 1 2
timestamp 1739975162
<< nwell >>
rect -38 262 774 582
<< pwell >>
rect 0 30 736 204
rect 0 28 644 30
rect 0 22 460 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 190 298 220 496
rect 286 298 316 496
rect 376 298 406 496
rect 472 298 502 496
rect 606 298 636 496
<< nmoslvt >>
rect 80 48 110 178
rect 190 48 220 178
rect 286 48 316 178
rect 376 48 406 178
rect 472 48 502 178
rect 606 48 636 178
<< ndiff >>
rect 27 94 80 178
rect 27 60 35 94
rect 69 60 80 94
rect 27 48 80 60
rect 110 150 190 178
rect 110 72 121 150
rect 155 72 190 150
rect 110 48 190 72
rect 220 48 286 178
rect 316 48 376 178
rect 406 94 472 178
rect 406 60 421 94
rect 455 60 472 94
rect 406 48 472 60
rect 502 170 606 178
rect 502 72 560 170
rect 594 72 606 170
rect 502 48 606 72
rect 636 136 708 178
rect 636 56 647 136
rect 681 56 708 136
rect 636 48 708 56
<< pdiff >>
rect 27 474 80 496
rect 27 314 35 474
rect 69 314 80 474
rect 27 298 80 314
rect 110 474 190 496
rect 110 400 130 474
rect 164 400 190 474
rect 110 298 190 400
rect 220 488 286 496
rect 220 454 231 488
rect 265 454 286 488
rect 220 298 286 454
rect 316 474 376 496
rect 316 400 327 474
rect 363 400 376 474
rect 316 298 376 400
rect 406 488 472 496
rect 406 318 417 488
rect 451 318 472 488
rect 406 298 472 318
rect 502 476 606 496
rect 502 306 560 476
rect 594 306 606 476
rect 502 298 606 306
rect 636 488 708 496
rect 636 340 647 488
rect 681 340 708 488
rect 636 298 708 340
<< ndiffc >>
rect 35 60 69 94
rect 121 72 155 150
rect 421 60 455 94
rect 560 72 594 170
rect 647 56 681 136
<< pdiffc >>
rect 35 314 69 474
rect 130 400 164 474
rect 231 454 265 488
rect 327 400 363 474
rect 417 318 451 488
rect 560 306 594 476
rect 647 340 681 488
<< poly >>
rect 80 496 110 522
rect 190 496 220 522
rect 286 496 316 522
rect 376 496 406 522
rect 472 496 502 522
rect 606 496 636 522
rect 80 268 110 298
rect 190 268 220 298
rect 286 268 316 298
rect 376 268 406 298
rect 472 268 502 298
rect 606 268 636 298
rect 80 250 142 268
rect 80 216 96 250
rect 130 216 142 250
rect 80 200 142 216
rect 184 250 238 268
rect 184 216 194 250
rect 228 216 238 250
rect 184 200 238 216
rect 280 250 334 268
rect 280 216 290 250
rect 324 216 334 250
rect 280 200 334 216
rect 376 250 430 268
rect 376 216 386 250
rect 420 216 430 250
rect 376 200 430 216
rect 472 250 636 268
rect 472 216 482 250
rect 516 216 636 250
rect 472 200 636 216
rect 80 178 110 200
rect 190 178 220 200
rect 286 178 316 200
rect 376 178 406 200
rect 472 178 502 200
rect 606 178 636 200
rect 80 22 110 48
rect 190 22 220 48
rect 286 22 316 48
rect 376 22 406 48
rect 472 22 502 48
rect 606 22 636 48
<< polycont >>
rect 96 216 130 250
rect 194 216 228 250
rect 290 216 324 250
rect 386 216 420 250
rect 482 216 516 250
<< locali >>
rect 0 561 736 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 526 736 527
rect 27 474 69 490
rect 27 314 35 474
rect 130 474 164 490
rect 231 488 265 526
rect 214 454 231 488
rect 265 454 282 488
rect 214 452 282 454
rect 327 474 363 490
rect 164 400 327 418
rect 130 384 363 400
rect 417 488 451 526
rect 27 298 69 314
rect 27 166 61 298
rect 104 268 142 350
rect 96 250 142 268
rect 130 216 142 250
rect 96 200 142 216
rect 178 250 228 350
rect 417 302 451 318
rect 560 476 594 492
rect 647 488 681 526
rect 647 324 681 340
rect 560 298 594 306
rect 178 216 194 250
rect 178 200 228 216
rect 262 250 334 268
rect 262 216 290 250
rect 324 216 334 250
rect 262 200 334 216
rect 376 250 430 268
rect 376 216 386 250
rect 420 216 430 250
rect 376 200 430 216
rect 472 250 526 268
rect 472 216 482 250
rect 516 216 526 250
rect 472 200 526 216
rect 27 150 155 166
rect 27 132 121 150
rect 19 94 85 98
rect 19 60 35 94
rect 69 60 85 94
rect 262 124 302 200
rect 472 162 508 200
rect 336 128 508 162
rect 560 178 624 298
rect 560 170 594 178
rect 336 90 370 128
rect 155 72 370 90
rect 35 21 69 60
rect 121 56 370 72
rect 405 60 421 94
rect 455 60 473 94
rect 421 21 455 60
rect 560 56 594 72
rect 647 136 681 152
rect 647 21 681 56
rect 0 17 736 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ao31_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 A
flabel locali s 272 221 306 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 289 238 289 238 0 FreeSans 200 0 0 0 B
flabel locali s 391 221 425 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 408 238 408 238 0 FreeSans 200 0 0 0 C
flabel locali s 102 221 136 255 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel locali s 119 238 119 238 0 FreeSans 200 0 0 0 D
flabel locali s 561 221 595 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 578 238 578 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__ao31_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 736 220
string MASKHINTS_NSDM 0 -38 736 209
string MASKHINTS_PSDM 0 273 736 582
<< end >>
