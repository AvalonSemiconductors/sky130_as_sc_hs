magic
tech sky130A
magscale 1 2
timestamp 1739438413
<< nwell >>
rect -38 262 774 582
<< pwell >>
rect 0 20 736 204
rect 26 -20 90 20
rect 486 -15 536 20
rect 486 -20 526 -15
<< pmos >>
rect 80 299 110 496
rect 166 299 196 496
rect 252 299 282 496
rect 338 299 368 496
rect 538 299 568 496
rect 624 299 654 496
<< nmoslvt >>
rect 80 49 110 178
rect 166 49 196 178
rect 252 49 282 178
rect 338 49 368 178
rect 538 49 568 178
rect 624 49 654 178
<< ndiff >>
rect 27 154 80 178
rect 27 62 35 154
rect 69 62 80 154
rect 27 49 80 62
rect 110 160 166 178
rect 110 72 121 160
rect 155 72 166 160
rect 110 49 166 72
rect 196 92 252 178
rect 196 58 207 92
rect 241 58 252 92
rect 196 49 252 58
rect 282 160 338 178
rect 282 72 293 160
rect 327 72 338 160
rect 282 49 338 72
rect 368 92 538 178
rect 368 58 380 92
rect 526 58 538 92
rect 368 49 538 58
rect 568 160 624 178
rect 568 72 579 160
rect 613 72 624 160
rect 568 49 624 72
rect 654 166 708 178
rect 654 62 665 166
rect 699 62 708 166
rect 654 49 708 62
<< pdiff >>
rect 27 474 80 496
rect 27 322 35 474
rect 69 322 80 474
rect 27 299 80 322
rect 110 488 166 496
rect 110 390 121 488
rect 155 390 166 488
rect 110 299 166 390
rect 196 474 252 496
rect 196 322 207 474
rect 241 322 252 474
rect 196 299 252 322
rect 282 406 338 496
rect 282 320 293 406
rect 327 320 338 406
rect 282 299 338 320
rect 368 474 430 496
rect 368 440 379 474
rect 413 440 430 474
rect 368 299 430 440
rect 484 474 538 496
rect 484 320 493 474
rect 527 320 538 474
rect 484 299 538 320
rect 568 406 624 496
rect 568 308 579 406
rect 613 308 624 406
rect 568 299 624 308
rect 654 474 708 496
rect 654 314 665 474
rect 699 314 708 474
rect 654 299 708 314
<< ndiffc >>
rect 35 62 69 154
rect 121 72 155 160
rect 207 58 241 92
rect 293 72 327 160
rect 380 58 526 92
rect 579 72 613 160
rect 665 62 699 166
<< pdiffc >>
rect 35 322 69 474
rect 121 390 155 488
rect 207 322 241 474
rect 293 320 327 406
rect 379 440 413 474
rect 493 320 527 474
rect 579 308 613 406
rect 665 314 699 474
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 538 496 568 522
rect 624 496 654 522
rect 80 268 110 299
rect 166 268 196 299
rect 252 268 282 299
rect 338 268 368 299
rect 62 252 196 268
rect 62 218 78 252
rect 180 218 196 252
rect 62 200 196 218
rect 238 252 370 268
rect 538 266 568 299
rect 624 266 654 299
rect 238 218 254 252
rect 358 218 370 252
rect 238 200 370 218
rect 442 252 656 266
rect 442 218 458 252
rect 510 218 656 252
rect 80 178 110 200
rect 166 178 196 200
rect 252 178 282 200
rect 338 178 368 200
rect 442 198 656 218
rect 538 178 568 198
rect 624 178 654 198
rect 80 23 110 49
rect 166 23 196 49
rect 252 23 282 49
rect 338 23 368 49
rect 538 23 568 49
rect 624 23 654 49
<< polycont >>
rect 78 218 180 252
rect 254 218 358 252
rect 458 218 510 252
<< locali >>
rect 0 561 736 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 526 736 527
rect 32 474 72 490
rect 32 322 35 474
rect 69 340 72 474
rect 114 488 162 526
rect 114 390 121 488
rect 155 390 162 488
rect 114 374 162 390
rect 204 474 416 490
rect 204 340 207 474
rect 69 322 207 340
rect 241 456 379 474
rect 241 322 244 456
rect 376 440 379 456
rect 413 440 416 474
rect 376 424 416 440
rect 490 474 704 490
rect 32 306 244 322
rect 290 406 330 422
rect 290 320 293 406
rect 327 390 330 406
rect 490 390 493 474
rect 327 356 493 390
rect 327 320 330 356
rect 290 302 330 320
rect 62 252 196 268
rect 62 218 78 252
rect 180 218 196 252
rect 62 212 196 218
rect 238 252 374 268
rect 238 218 254 252
rect 358 218 374 252
rect 422 262 456 322
rect 490 320 493 356
rect 527 456 665 474
rect 527 320 530 456
rect 490 302 530 320
rect 574 406 616 422
rect 574 308 579 406
rect 613 308 616 406
rect 574 292 616 308
rect 664 314 665 456
rect 699 314 704 474
rect 664 298 704 314
rect 422 252 526 262
rect 422 218 458 252
rect 510 218 526 252
rect 238 212 374 218
rect 574 176 620 292
rect 121 174 620 176
rect 35 154 69 170
rect 35 21 69 62
rect 121 160 613 174
rect 155 142 293 160
rect 121 56 155 72
rect 207 92 241 108
rect 207 21 241 58
rect 327 142 579 160
rect 293 56 327 72
rect 380 92 530 108
rect 526 58 530 92
rect 380 21 530 58
rect 579 56 613 72
rect 665 166 699 182
rect 665 21 699 62
rect 0 17 736 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor3_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 A
flabel locali 255 221 289 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 272 238 272 238 0 FreeSans 200 0 0 0 B
flabel locali 459 221 493 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel polycont 476 238 476 238 0 FreeSans 200 0 0 0 C
flabel locali 578 221 612 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali 595 238 595 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor3_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 736 216
string MASKHINTS_NSDM 0 -38 736 204
string MASKHINTS_PSDM 0 272 736 582
<< end >>
