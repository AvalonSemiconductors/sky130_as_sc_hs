magic
tech sky130A
magscale 1 2
timestamp 1733957473
<< nwell >>
rect -38 262 314 582
<< pwell >>
rect 0 -18 276 204
<< nmoslvt >>
rect 80 50 110 183
rect 166 50 196 183
<< pmos >>
rect 80 314 110 497
rect 166 314 196 497
<< ndiff >>
rect 27 156 80 183
rect 27 74 35 156
rect 69 74 80 156
rect 27 50 80 74
rect 110 158 166 183
rect 110 76 121 158
rect 155 76 166 158
rect 110 50 166 76
rect 196 167 249 183
rect 196 94 207 167
rect 241 94 249 167
rect 196 50 249 94
<< pdiff >>
rect 27 485 80 497
rect 27 348 35 485
rect 69 348 80 485
rect 27 314 80 348
rect 110 314 166 497
rect 196 476 249 497
rect 196 346 207 476
rect 241 346 249 476
rect 196 314 249 346
<< ndiffc >>
rect 35 74 69 156
rect 121 76 155 158
rect 207 94 241 167
<< pdiffc >>
rect 35 348 69 485
rect 207 346 241 476
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 80 282 110 314
rect 25 266 110 282
rect 25 232 35 266
rect 69 232 110 266
rect 25 216 110 232
rect 80 183 110 216
rect 166 284 196 314
rect 166 267 249 284
rect 166 233 205 267
rect 239 233 249 267
rect 166 217 249 233
rect 166 183 196 217
rect 80 24 110 50
rect 166 24 196 50
<< polycont >>
rect 35 232 69 266
rect 205 233 239 267
<< locali >>
rect 0 561 276 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 526 276 527
rect 35 485 69 526
rect 207 476 241 492
rect 35 322 69 348
rect 121 346 207 356
rect 121 322 241 346
rect 33 266 87 284
rect 33 232 35 266
rect 69 232 87 266
rect 33 216 87 232
rect 121 176 155 322
rect 189 267 241 286
rect 189 233 205 267
rect 239 233 241 267
rect 189 217 241 233
rect 35 156 69 172
rect 115 158 155 176
rect 115 134 121 158
rect 35 21 69 74
rect 121 60 155 76
rect 207 167 241 183
rect 207 21 241 94
rect 0 17 276 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor2_1
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 276 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 276 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 204 238 238 272 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali s 221 255 221 255 0 FreeSans 200 0 0 0 B
flabel locali s 119 136 153 170 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel ndiffc 136 153 136 153 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor2_1.mag
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 6.900 0.000 
<< end >>
