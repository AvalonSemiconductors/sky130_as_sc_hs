magic
tech sky130A
magscale 1 2
timestamp 1740276425
<< nwell >>
rect -38 262 682 582
<< pwell >>
rect 10 48 644 204
rect 26 44 320 48
rect 26 26 90 44
rect 372 30 644 48
rect 26 22 110 26
rect 26 -20 90 22
<< pmos >>
rect 80 314 110 496
rect 166 314 196 496
rect 264 314 294 496
rect 350 314 380 496
rect 436 314 466 496
rect 522 314 552 496
<< nmoslvt >>
rect 80 48 110 184
rect 166 48 196 184
rect 264 48 294 184
rect 350 48 380 184
rect 436 48 466 184
rect 522 48 552 184
<< ndiff >>
rect 27 166 80 184
rect 27 72 35 166
rect 69 72 80 166
rect 27 48 80 72
rect 110 48 166 184
rect 196 156 264 184
rect 196 72 207 156
rect 241 72 264 156
rect 196 48 264 72
rect 294 166 350 184
rect 294 72 305 166
rect 339 72 350 166
rect 294 48 350 72
rect 380 102 436 184
rect 380 61 391 102
rect 425 61 436 102
rect 380 48 436 61
rect 466 176 522 184
rect 466 72 477 176
rect 511 72 522 176
rect 466 48 522 72
rect 552 168 617 184
rect 552 56 563 168
rect 597 56 617 168
rect 552 48 617 56
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 314 80 336
rect 110 476 166 496
rect 110 348 121 476
rect 155 348 166 476
rect 110 314 166 348
rect 196 488 264 496
rect 196 406 207 488
rect 241 406 264 488
rect 196 314 264 406
rect 294 474 350 496
rect 294 406 305 474
rect 339 406 350 474
rect 294 314 350 406
rect 380 484 436 496
rect 380 450 391 484
rect 425 450 436 484
rect 380 314 436 450
rect 466 474 522 496
rect 466 322 477 474
rect 511 322 522 474
rect 466 314 522 322
rect 552 488 617 496
rect 552 330 563 488
rect 597 330 617 488
rect 552 314 617 330
<< ndiffc >>
rect 35 72 69 166
rect 207 72 241 156
rect 305 72 339 166
rect 391 61 425 102
rect 477 72 511 176
rect 563 56 597 168
<< pdiffc >>
rect 35 336 69 476
rect 121 348 155 476
rect 207 406 241 488
rect 305 406 339 474
rect 391 450 425 484
rect 477 322 511 474
rect 563 330 597 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 264 496 294 522
rect 350 496 380 522
rect 436 496 466 522
rect 522 496 552 522
rect 80 284 110 314
rect 30 266 110 284
rect 30 232 42 266
rect 76 232 110 266
rect 30 216 110 232
rect 80 184 110 216
rect 166 284 196 314
rect 264 288 294 314
rect 350 288 380 314
rect 436 288 466 314
rect 522 288 552 314
rect 166 266 222 284
rect 166 232 178 266
rect 212 232 222 266
rect 166 212 222 232
rect 264 266 552 288
rect 264 232 274 266
rect 308 232 552 266
rect 264 216 552 232
rect 166 184 196 212
rect 264 184 294 216
rect 350 184 380 216
rect 436 184 466 216
rect 522 184 552 216
rect 80 22 110 48
rect 166 22 196 48
rect 264 22 294 48
rect 350 22 380 48
rect 436 22 466 48
rect 522 22 552 48
<< polycont >>
rect 42 232 76 266
rect 178 232 212 266
rect 274 232 308 266
<< locali >>
rect 0 561 644 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 526 644 527
rect 35 476 69 526
rect 121 476 155 492
rect 35 320 69 336
rect 110 348 121 362
rect 207 488 241 526
rect 207 390 241 406
rect 303 474 340 490
rect 303 406 305 474
rect 339 416 340 474
rect 374 484 442 526
rect 374 450 391 484
rect 425 450 442 484
rect 477 474 511 490
rect 339 406 400 416
rect 303 390 400 406
rect 312 382 400 390
rect 155 348 290 356
rect 110 320 290 348
rect 30 266 76 286
rect 30 232 42 266
rect 30 216 76 232
rect 110 182 144 320
rect 256 288 290 320
rect 342 292 400 382
rect 477 292 511 322
rect 563 488 597 526
rect 563 314 597 330
rect 178 266 222 282
rect 212 232 222 266
rect 178 214 222 232
rect 256 266 308 288
rect 256 232 274 266
rect 256 216 308 232
rect 342 220 511 292
rect 342 182 400 220
rect 34 166 144 182
rect 34 148 35 166
rect 69 148 144 166
rect 207 156 241 176
rect 35 56 69 72
rect 207 21 241 72
rect 303 166 400 182
rect 303 72 305 166
rect 339 154 400 166
rect 477 176 511 220
rect 339 148 374 154
rect 303 56 339 72
rect 391 102 425 118
rect 391 21 425 61
rect 477 56 511 72
rect 563 168 597 184
rect 563 21 597 56
rect 0 17 644 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
flabel locali 187 221 221 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 204 238 204 238 0 FreeSans 200 0 0 0 B
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__and2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 644 220
string MASKHINTS_NSDM 0 -38 644 209
string MASKHINTS_PSDM 0 289 644 582
<< end >>
