magic
tech sky130A
magscale 1 2
timestamp 1739438880
<< nwell >>
rect -38 262 866 582
<< pwell >>
rect 0 28 828 204
rect 0 22 736 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 152 298 182 496
rect 238 298 268 496
rect 310 298 340 496
rect 396 298 426 496
rect 468 298 498 496
rect 576 298 606 496
rect 662 298 692 496
<< nmoslvt >>
rect 80 49 110 178
rect 152 49 182 178
rect 238 49 268 178
rect 310 49 340 178
rect 396 49 426 178
rect 468 49 498 178
rect 576 49 606 178
rect 662 49 692 178
<< ndiff >>
rect 27 164 80 178
rect 27 72 35 164
rect 69 72 80 164
rect 27 49 80 72
rect 110 49 152 178
rect 182 96 238 178
rect 182 58 193 96
rect 227 58 238 96
rect 182 49 238 58
rect 268 49 310 178
rect 340 170 396 178
rect 340 72 351 170
rect 385 72 396 170
rect 340 49 396 72
rect 426 49 468 178
rect 498 96 576 178
rect 498 58 520 96
rect 554 58 576 96
rect 498 49 576 58
rect 606 110 662 178
rect 606 76 617 110
rect 651 76 662 110
rect 606 49 662 76
rect 692 164 801 178
rect 692 58 744 164
rect 778 58 801 164
rect 692 49 801 58
<< pdiff >>
rect 27 476 80 496
rect 27 386 35 476
rect 69 386 80 476
rect 27 298 80 386
rect 110 298 152 496
rect 182 488 238 496
rect 182 454 193 488
rect 227 454 238 488
rect 182 298 238 454
rect 268 298 310 496
rect 340 476 396 496
rect 340 370 351 476
rect 385 370 396 476
rect 340 298 396 370
rect 426 298 468 496
rect 498 488 576 496
rect 498 454 509 488
rect 543 454 576 488
rect 498 298 576 454
rect 606 464 662 496
rect 606 430 617 464
rect 651 430 662 464
rect 606 298 662 430
rect 692 488 801 496
rect 692 306 744 488
rect 778 306 801 488
rect 692 298 801 306
<< ndiffc >>
rect 35 72 69 164
rect 193 58 227 96
rect 351 72 385 170
rect 520 58 554 96
rect 617 76 651 110
rect 744 58 778 164
<< pdiffc >>
rect 35 386 69 476
rect 193 454 227 488
rect 351 370 385 476
rect 509 454 543 488
rect 617 430 651 464
rect 744 306 778 488
<< poly >>
rect 80 496 110 522
rect 152 496 182 522
rect 238 496 268 522
rect 310 496 340 522
rect 396 496 426 522
rect 468 496 498 522
rect 576 496 606 522
rect 662 496 692 522
rect 80 266 110 298
rect 44 250 110 266
rect 44 216 60 250
rect 94 216 110 250
rect 44 204 110 216
rect 80 178 110 204
rect 152 266 182 298
rect 238 266 268 298
rect 152 250 268 266
rect 152 216 168 250
rect 252 216 268 250
rect 152 204 268 216
rect 152 178 182 204
rect 238 178 268 204
rect 310 266 340 298
rect 396 266 426 298
rect 310 250 426 266
rect 310 216 326 250
rect 410 216 426 250
rect 310 204 426 216
rect 310 178 340 204
rect 396 178 426 204
rect 468 266 498 298
rect 576 266 606 298
rect 662 266 692 298
rect 468 250 534 266
rect 468 216 484 250
rect 518 216 534 250
rect 468 204 534 216
rect 576 250 692 266
rect 576 216 592 250
rect 626 216 692 250
rect 576 204 692 216
rect 468 178 498 204
rect 576 178 606 204
rect 662 178 692 204
rect 80 23 110 49
rect 152 23 182 49
rect 238 23 268 49
rect 310 23 340 49
rect 396 23 426 49
rect 468 23 498 49
rect 576 23 606 49
rect 662 23 692 49
<< polycont >>
rect 60 216 94 250
rect 168 216 252 250
rect 326 216 410 250
rect 484 216 518 250
rect 592 216 626 250
<< locali >>
rect 0 561 828 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 526 828 527
rect 34 476 70 492
rect 34 386 35 476
rect 69 404 70 476
rect 193 488 227 526
rect 193 438 227 454
rect 350 476 386 492
rect 350 404 351 476
rect 69 386 351 404
rect 34 370 351 386
rect 385 404 386 476
rect 509 488 543 526
rect 744 488 778 526
rect 509 438 543 454
rect 617 464 651 488
rect 651 430 710 448
rect 617 414 710 430
rect 385 372 570 404
rect 385 370 602 372
rect 536 338 602 370
rect 70 300 502 334
rect 70 266 110 300
rect 468 266 502 300
rect 568 266 602 338
rect 44 250 110 266
rect 44 216 60 250
rect 94 216 110 250
rect 44 214 110 216
rect 152 250 268 266
rect 152 216 168 250
rect 252 216 268 250
rect 152 214 268 216
rect 310 250 432 266
rect 310 216 326 250
rect 410 216 432 250
rect 310 214 432 216
rect 468 250 534 266
rect 468 216 484 250
rect 518 216 534 250
rect 468 214 534 216
rect 568 250 642 266
rect 568 216 592 250
rect 626 216 642 250
rect 568 214 642 216
rect 676 262 710 414
rect 744 290 778 306
rect 568 180 602 214
rect 35 170 602 180
rect 35 164 351 170
rect 69 146 351 164
rect 35 56 69 72
rect 193 96 227 112
rect 193 21 227 58
rect 385 146 602 170
rect 676 208 724 262
rect 351 56 385 72
rect 520 96 554 112
rect 676 110 710 208
rect 520 21 554 58
rect 600 76 617 110
rect 651 76 710 110
rect 744 164 778 180
rect 600 56 666 76
rect 744 21 778 58
rect 0 17 828 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel comment s 0 0 0 0 4 maj3_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 170 221 204 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 51 221 85 255 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 68 238 68 238 0 FreeSans 200 0 0 0 A
flabel locali 323 221 357 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali 340 238 340 238 0 FreeSans 200 0 0 0 C
flabel locali 680 221 714 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali 697 238 697 238 0 FreeSans 200 0 0 0 Y
flabel polycont 187 238 187 238 0 FreeSans 200 0 0 0 B
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__maj3_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 828 214
string MASKHINTS_NSDM 0 -38 828 204
string MASKHINTS_PSDM 0 272 828 582
<< end >>
