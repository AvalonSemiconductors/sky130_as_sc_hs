magic
tech sky130A
magscale 1 2
timestamp 1739569896
<< nwell >>
rect -38 262 1786 582
<< pwell >>
rect 18 48 1742 204
rect 22 44 1608 48
rect 22 -15 82 44
rect 22 -20 64 -15
<< pmos >>
rect 83 301 113 496
rect 170 301 200 496
rect 368 372 398 496
rect 466 401 496 496
rect 584 401 614 496
rect 754 393 784 496
rect 854 393 884 496
rect 962 393 992 496
rect 1076 385 1106 496
rect 1250 385 1280 496
rect 1352 385 1382 496
rect 1542 298 1572 496
rect 1628 298 1658 496
<< nmoslvt >>
rect 83 48 113 182
rect 170 48 200 182
rect 368 49 398 140
rect 468 49 498 138
rect 654 49 684 138
rect 754 49 784 144
rect 854 49 884 148
rect 964 49 994 138
rect 1150 49 1180 138
rect 1250 49 1280 148
rect 1352 49 1382 148
rect 1542 48 1572 178
rect 1628 48 1658 178
<< ndiff >>
rect 30 128 83 182
rect 30 72 38 128
rect 72 72 83 128
rect 30 48 83 72
rect 113 91 170 182
rect 113 57 124 91
rect 158 57 170 91
rect 113 48 170 57
rect 200 106 258 182
rect 200 72 212 106
rect 246 72 258 106
rect 200 48 258 72
rect 312 122 368 140
rect 312 64 322 122
rect 356 64 368 122
rect 312 49 368 64
rect 398 138 448 140
rect 804 144 854 148
rect 704 138 754 144
rect 398 130 468 138
rect 398 72 416 130
rect 450 72 468 130
rect 398 49 468 72
rect 498 120 654 138
rect 498 86 526 120
rect 560 86 654 120
rect 498 49 654 86
rect 684 49 754 138
rect 784 114 854 144
rect 784 60 806 114
rect 840 60 854 114
rect 784 49 854 60
rect 884 138 934 148
rect 1489 150 1542 178
rect 1200 138 1250 148
rect 884 130 964 138
rect 884 74 910 130
rect 944 74 964 130
rect 884 49 964 74
rect 994 120 1150 138
rect 994 86 1022 120
rect 1056 86 1150 120
rect 994 49 1150 86
rect 1180 49 1250 138
rect 1280 114 1352 148
rect 1280 60 1304 114
rect 1338 60 1352 114
rect 1280 49 1352 60
rect 1382 126 1435 148
rect 1382 72 1393 126
rect 1427 72 1435 126
rect 1382 49 1435 72
rect 1489 68 1497 150
rect 1531 68 1542 150
rect 1489 48 1542 68
rect 1572 170 1628 178
rect 1572 76 1583 170
rect 1617 76 1628 170
rect 1572 48 1628 76
rect 1658 166 1711 178
rect 1658 68 1669 166
rect 1703 68 1711 166
rect 1658 48 1711 68
<< pdiff >>
rect 28 470 83 496
rect 28 378 38 470
rect 72 378 83 470
rect 28 301 83 378
rect 113 484 170 496
rect 113 434 124 484
rect 158 434 170 484
rect 113 301 170 434
rect 200 470 258 496
rect 200 374 212 470
rect 246 374 258 470
rect 200 301 258 374
rect 312 484 368 496
rect 312 432 322 484
rect 356 432 368 484
rect 312 372 368 432
rect 398 472 466 496
rect 398 432 416 472
rect 450 432 466 472
rect 398 401 466 432
rect 496 476 584 496
rect 496 442 526 476
rect 560 442 584 476
rect 496 401 584 442
rect 614 401 754 496
rect 398 372 448 401
rect 680 393 754 401
rect 784 488 854 496
rect 784 432 798 488
rect 832 432 854 488
rect 784 393 854 432
rect 884 474 962 496
rect 884 420 910 474
rect 944 420 962 474
rect 884 393 962 420
rect 992 476 1076 496
rect 992 442 1022 476
rect 1056 442 1076 476
rect 992 393 1076 442
rect 1026 385 1076 393
rect 1106 385 1250 496
rect 1280 488 1352 496
rect 1280 432 1302 488
rect 1336 432 1352 488
rect 1280 385 1352 432
rect 1382 476 1435 496
rect 1382 422 1393 476
rect 1427 422 1435 476
rect 1382 385 1435 422
rect 1489 478 1542 496
rect 1489 388 1497 478
rect 1531 388 1542 478
rect 1489 298 1542 388
rect 1572 468 1628 496
rect 1572 306 1583 468
rect 1617 306 1628 468
rect 1572 298 1628 306
rect 1658 480 1711 496
rect 1658 310 1669 480
rect 1703 310 1711 480
rect 1658 298 1711 310
<< ndiffc >>
rect 38 72 72 128
rect 124 57 158 91
rect 212 72 246 106
rect 322 64 356 122
rect 416 72 450 130
rect 526 86 560 120
rect 806 60 840 114
rect 910 74 944 130
rect 1022 86 1056 120
rect 1304 60 1338 114
rect 1393 72 1427 126
rect 1497 68 1531 150
rect 1583 76 1617 170
rect 1669 68 1703 166
<< pdiffc >>
rect 38 378 72 470
rect 124 434 158 484
rect 212 374 246 470
rect 322 432 356 484
rect 416 432 450 472
rect 526 442 560 476
rect 798 432 832 488
rect 910 420 944 474
rect 1022 442 1056 476
rect 1302 432 1336 488
rect 1393 422 1427 476
rect 1497 388 1531 478
rect 1583 306 1617 468
rect 1669 310 1703 480
<< poly >>
rect 83 496 113 522
rect 170 496 200 522
rect 368 496 398 522
rect 466 496 496 522
rect 584 496 614 522
rect 754 496 784 522
rect 854 496 884 522
rect 962 496 992 522
rect 1076 496 1106 522
rect 1250 496 1280 522
rect 1352 496 1382 522
rect 1542 496 1572 522
rect 1628 496 1658 522
rect 83 267 113 301
rect 38 254 113 267
rect 38 220 54 254
rect 88 220 113 254
rect 38 208 113 220
rect 83 182 113 208
rect 170 270 200 301
rect 368 300 398 372
rect 466 364 496 401
rect 466 354 542 364
rect 466 320 492 354
rect 526 320 542 354
rect 466 310 542 320
rect 316 290 398 300
rect 170 254 228 270
rect 170 220 180 254
rect 214 220 228 254
rect 316 256 332 290
rect 366 256 398 290
rect 584 276 614 401
rect 574 268 614 276
rect 316 246 398 256
rect 170 204 228 220
rect 170 182 200 204
rect 368 140 398 246
rect 462 248 614 268
rect 462 214 482 248
rect 520 246 614 248
rect 754 262 784 393
rect 854 356 884 393
rect 826 346 888 356
rect 826 312 842 346
rect 876 312 888 346
rect 826 302 888 312
rect 962 348 992 393
rect 962 338 1034 348
rect 962 304 980 338
rect 1018 304 1034 338
rect 754 246 812 262
rect 520 238 596 246
rect 520 214 536 238
rect 462 204 536 214
rect 654 216 712 232
rect 468 138 498 204
rect 654 182 664 216
rect 702 182 712 216
rect 654 166 712 182
rect 754 212 764 246
rect 802 212 812 246
rect 754 196 812 212
rect 654 138 684 166
rect 754 144 784 196
rect 854 148 884 302
rect 962 294 1034 304
rect 1076 252 1106 385
rect 964 238 1106 252
rect 964 204 984 238
rect 1022 222 1106 238
rect 1150 232 1208 248
rect 1022 204 1038 222
rect 964 194 1038 204
rect 1150 198 1160 232
rect 1198 198 1208 232
rect 964 138 994 194
rect 1150 182 1208 198
rect 1250 246 1280 385
rect 1352 342 1382 385
rect 1322 332 1384 342
rect 1322 298 1338 332
rect 1372 298 1384 332
rect 1322 288 1384 298
rect 1250 230 1308 246
rect 1250 196 1260 230
rect 1298 196 1308 230
rect 1150 138 1180 182
rect 1250 180 1308 196
rect 1250 148 1280 180
rect 1352 148 1382 288
rect 1542 270 1572 298
rect 1628 270 1658 298
rect 1444 250 1658 270
rect 1444 216 1460 250
rect 1494 216 1658 250
rect 1444 206 1658 216
rect 1444 200 1572 206
rect 1542 178 1572 200
rect 1628 178 1658 206
rect 83 22 113 48
rect 170 22 200 48
rect 368 23 398 49
rect 468 23 498 49
rect 654 23 684 49
rect 754 23 784 49
rect 854 23 884 49
rect 964 23 994 49
rect 1150 23 1180 49
rect 1250 23 1280 49
rect 1352 23 1382 49
rect 1542 22 1572 48
rect 1628 22 1658 48
<< polycont >>
rect 54 220 88 254
rect 492 320 526 354
rect 180 220 214 254
rect 332 256 366 290
rect 482 214 520 248
rect 842 312 876 346
rect 980 304 1018 338
rect 664 182 702 216
rect 764 212 802 246
rect 984 204 1022 238
rect 1160 198 1198 232
rect 1338 298 1372 332
rect 1260 196 1298 230
rect 1460 216 1494 250
<< locali >>
rect 0 561 1748 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 526 1748 527
rect 38 470 72 488
rect 124 484 158 526
rect 124 418 158 434
rect 212 470 246 488
rect 72 378 156 384
rect 38 350 156 378
rect 322 484 356 526
rect 322 414 356 432
rect 416 472 450 490
rect 798 488 832 526
rect 510 442 526 476
rect 416 414 450 432
rect 246 374 282 384
rect 212 360 282 374
rect 212 350 248 360
rect 28 254 88 316
rect 28 220 54 254
rect 28 196 88 220
rect 122 270 156 350
rect 242 326 248 350
rect 410 344 450 414
rect 484 368 526 370
rect 242 318 282 326
rect 122 254 214 270
rect 122 220 180 254
rect 122 204 214 220
rect 122 162 156 204
rect 38 128 122 162
rect 248 122 282 318
rect 316 290 376 336
rect 316 256 332 290
rect 366 256 376 290
rect 316 184 376 256
rect 410 176 444 344
rect 484 334 488 368
rect 484 320 492 334
rect 484 304 526 320
rect 560 356 594 476
rect 798 416 832 432
rect 910 474 944 490
rect 1302 488 1336 526
rect 1006 442 1022 476
rect 834 356 876 362
rect 560 346 876 356
rect 560 322 842 346
rect 478 260 520 264
rect 478 248 486 260
rect 478 214 482 248
rect 478 198 520 214
rect 212 106 282 122
rect 38 56 72 72
rect 108 91 174 94
rect 108 57 124 91
rect 158 57 174 91
rect 108 56 174 57
rect 246 72 282 106
rect 212 56 282 72
rect 322 122 356 150
rect 410 138 450 176
rect 560 164 594 322
rect 834 312 842 322
rect 834 296 876 312
rect 760 246 802 262
rect 910 246 944 420
rect 978 362 1020 366
rect 978 304 980 362
rect 1018 304 1020 362
rect 978 288 1020 304
rect 1056 358 1090 476
rect 1302 416 1336 432
rect 1388 476 1440 492
rect 1388 422 1393 476
rect 1427 422 1440 476
rect 1388 406 1440 422
rect 1056 332 1372 358
rect 1056 324 1338 332
rect 660 216 702 232
rect 660 180 664 216
rect 760 212 764 246
rect 802 212 944 246
rect 760 196 802 212
rect 660 166 702 180
rect 124 21 158 56
rect 322 21 356 64
rect 416 130 450 138
rect 542 130 594 164
rect 910 130 944 212
rect 980 250 1022 254
rect 980 204 984 250
rect 980 188 1022 204
rect 1056 130 1090 324
rect 1334 298 1338 324
rect 1334 282 1372 298
rect 1406 270 1440 406
rect 1497 478 1531 526
rect 1497 372 1531 388
rect 1578 468 1622 484
rect 1578 338 1583 468
rect 1538 306 1583 338
rect 1617 306 1622 468
rect 1406 250 1504 270
rect 1158 232 1200 248
rect 1158 182 1160 232
rect 1198 182 1200 232
rect 1158 176 1200 182
rect 1256 246 1298 248
rect 1406 246 1460 250
rect 1256 230 1460 246
rect 1256 196 1260 230
rect 1298 216 1460 230
rect 1494 216 1504 250
rect 1538 230 1622 306
rect 1669 480 1703 526
rect 1669 294 1703 310
rect 1298 212 1504 216
rect 1256 180 1298 196
rect 1406 200 1504 212
rect 1406 158 1440 200
rect 1578 170 1622 230
rect 1391 134 1440 158
rect 1497 150 1531 166
rect 542 120 576 130
rect 510 86 526 120
rect 560 86 576 120
rect 806 114 840 130
rect 416 56 450 72
rect 806 21 840 60
rect 1038 120 1090 130
rect 1006 86 1022 120
rect 1056 86 1090 120
rect 1304 114 1338 130
rect 910 58 944 74
rect 1304 21 1338 60
rect 1391 126 1432 134
rect 1391 72 1393 126
rect 1427 72 1432 126
rect 1391 56 1432 72
rect 1497 21 1531 68
rect 1578 76 1583 170
rect 1617 76 1622 170
rect 1578 60 1622 76
rect 1669 166 1703 182
rect 1669 21 1703 68
rect 0 17 1748 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 248 326 282 360
rect 122 128 156 162
rect 488 354 526 368
rect 488 334 492 354
rect 492 334 526 354
rect 486 248 520 260
rect 486 226 520 248
rect 980 338 1018 362
rect 980 328 1018 338
rect 664 182 702 216
rect 664 180 702 182
rect 984 238 1022 250
rect 984 212 1022 238
rect 1160 198 1198 216
rect 1160 182 1198 198
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 482 368 532 376
rect 234 360 488 368
rect 234 326 248 360
rect 282 334 488 360
rect 526 334 878 368
rect 282 326 294 334
rect 482 328 532 334
rect 234 318 294 326
rect 474 260 532 268
rect 474 226 486 260
rect 520 226 532 260
rect 660 238 694 334
rect 842 264 878 334
rect 968 362 1198 368
rect 968 328 980 362
rect 1018 328 1198 362
rect 968 322 1198 328
rect 972 264 1034 266
rect 842 250 1034 264
rect 474 220 532 226
rect 500 218 532 220
rect 110 162 184 168
rect 110 128 122 162
rect 156 128 184 162
rect 110 126 184 128
rect 500 128 528 218
rect 658 216 708 238
rect 842 230 984 250
rect 658 180 664 216
rect 702 180 708 216
rect 972 212 984 230
rect 1022 212 1034 250
rect 1154 238 1198 322
rect 972 206 1034 212
rect 1152 216 1206 238
rect 658 164 708 180
rect 1152 182 1160 216
rect 1198 182 1206 216
rect 1152 164 1206 182
rect 1172 128 1200 164
rect 500 126 1200 128
rect 110 116 1200 126
rect 150 98 1200 116
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxtp_2
flabel locali s 29 272 63 306 0 FreeSans 400 0 0 0 CLK
port 5 nsew clock input
flabel locali s 46 289 46 289 0 FreeSans 400 0 0 0 CLK
flabel locali s 329 238 363 272 0 FreeSans 200 0 0 0 D
port 7 nsew signal input
flabel locali s 346 255 346 255 0 FreeSans 200 0 0 0 D
flabel locali s 1569 272 1603 306 0 FreeSans 200 0 0 0 Q
port 6 nsew signal output
flabel locali s 1586 289 1586 289 0 FreeSans 200 0 0 0 Q
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel metal1 s 0 -48 1748 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__dfxtp_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1748 218
string MASKHINTS_NSDM 0 -38 1748 207
string MASKHINTS_PSDM 0 272 1748 582
<< end >>
