magic
tech sky130A
magscale 1 2
timestamp 1739658706
<< nwell >>
rect -38 262 1510 582
<< pwell >>
rect 456 206 1336 220
rect 20 44 1424 204
rect 20 -15 82 44
rect 20 -20 74 -15
<< pmos >>
rect 81 312 111 496
rect 168 312 198 496
rect 256 312 286 496
rect 344 312 374 496
rect 432 312 462 496
rect 524 312 554 496
rect 612 312 642 496
rect 700 312 730 496
rect 788 312 818 496
rect 876 312 906 496
rect 964 312 994 496
rect 1052 312 1082 496
rect 1140 312 1170 496
rect 1230 312 1260 496
rect 1318 312 1348 496
<< nmoslvt >>
rect 81 48 111 179
rect 168 48 198 179
rect 256 48 286 179
rect 344 48 374 179
rect 432 48 462 179
rect 524 48 554 179
rect 612 48 642 179
rect 700 48 730 179
rect 788 48 818 179
rect 876 48 906 179
rect 964 48 994 179
rect 1052 48 1082 179
rect 1140 48 1170 179
rect 1230 48 1260 179
rect 1318 48 1348 179
<< ndiff >>
rect 28 132 81 179
rect 28 64 36 132
rect 70 64 81 132
rect 28 48 81 64
rect 111 150 168 179
rect 111 72 122 150
rect 156 72 168 150
rect 111 48 168 72
rect 198 98 256 179
rect 198 64 210 98
rect 244 64 256 98
rect 198 48 256 64
rect 286 150 344 179
rect 286 72 298 150
rect 332 72 344 150
rect 286 48 344 72
rect 374 98 432 179
rect 374 64 386 98
rect 420 64 432 98
rect 374 48 432 64
rect 462 150 524 179
rect 462 72 478 150
rect 512 72 524 150
rect 462 48 524 72
rect 554 99 612 179
rect 554 64 566 99
rect 600 64 612 99
rect 554 48 612 64
rect 642 150 700 179
rect 642 72 654 150
rect 688 72 700 150
rect 642 48 700 72
rect 730 95 788 179
rect 730 60 742 95
rect 776 60 788 95
rect 730 48 788 60
rect 818 150 876 179
rect 818 72 830 150
rect 864 72 876 150
rect 818 48 876 72
rect 906 95 964 179
rect 906 60 918 95
rect 952 60 964 95
rect 906 48 964 60
rect 994 150 1052 179
rect 994 72 1006 150
rect 1040 72 1052 150
rect 994 48 1052 72
rect 1082 99 1140 179
rect 1082 58 1094 99
rect 1128 58 1140 99
rect 1082 48 1140 58
rect 1170 150 1230 179
rect 1170 72 1182 150
rect 1216 72 1230 150
rect 1170 48 1230 72
rect 1260 99 1318 179
rect 1260 58 1272 99
rect 1306 58 1318 99
rect 1260 48 1318 58
rect 1348 150 1406 179
rect 1348 72 1360 150
rect 1394 72 1406 150
rect 1348 48 1406 72
<< pdiff >>
rect 28 480 81 496
rect 28 394 36 480
rect 70 394 81 480
rect 28 312 81 394
rect 111 476 168 496
rect 111 360 122 476
rect 156 360 168 476
rect 111 312 168 360
rect 198 482 256 496
rect 198 407 210 482
rect 244 407 256 482
rect 198 312 256 407
rect 286 476 344 496
rect 286 360 298 476
rect 332 360 344 476
rect 286 312 344 360
rect 374 484 432 496
rect 374 408 386 484
rect 420 408 432 484
rect 374 312 432 408
rect 462 476 524 496
rect 462 322 478 476
rect 512 322 524 476
rect 462 312 524 322
rect 554 484 612 496
rect 554 409 566 484
rect 600 409 612 484
rect 554 312 612 409
rect 642 476 700 496
rect 642 320 654 476
rect 688 320 700 476
rect 642 312 700 320
rect 730 484 788 496
rect 730 409 742 484
rect 776 409 788 484
rect 730 312 788 409
rect 818 476 876 496
rect 818 320 830 476
rect 864 320 876 476
rect 818 312 876 320
rect 906 484 964 496
rect 906 409 918 484
rect 952 409 964 484
rect 906 312 964 409
rect 994 476 1052 496
rect 994 320 1006 476
rect 1040 320 1052 476
rect 994 312 1052 320
rect 1082 484 1140 496
rect 1082 409 1094 484
rect 1128 409 1140 484
rect 1082 312 1140 409
rect 1170 476 1230 496
rect 1170 320 1184 476
rect 1218 320 1230 476
rect 1170 312 1230 320
rect 1260 484 1318 496
rect 1260 409 1272 484
rect 1306 409 1318 484
rect 1260 312 1318 409
rect 1348 476 1406 496
rect 1348 320 1360 476
rect 1394 320 1406 476
rect 1348 312 1406 320
<< ndiffc >>
rect 36 64 70 132
rect 122 72 156 150
rect 210 64 244 98
rect 298 72 332 150
rect 386 64 420 98
rect 478 72 512 150
rect 566 64 600 99
rect 654 72 688 150
rect 742 60 776 95
rect 830 72 864 150
rect 918 60 952 95
rect 1006 72 1040 150
rect 1094 58 1128 99
rect 1182 72 1216 150
rect 1272 58 1306 99
rect 1360 72 1394 150
<< pdiffc >>
rect 36 394 70 480
rect 122 360 156 476
rect 210 407 244 482
rect 298 360 332 476
rect 386 408 420 484
rect 478 322 512 476
rect 566 409 600 484
rect 654 320 688 476
rect 742 409 776 484
rect 830 320 864 476
rect 918 409 952 484
rect 1006 320 1040 476
rect 1094 409 1128 484
rect 1184 320 1218 476
rect 1272 409 1306 484
rect 1360 320 1394 476
<< poly >>
rect 81 496 111 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 524 496 554 522
rect 612 496 642 522
rect 700 496 730 522
rect 788 496 818 522
rect 876 496 906 522
rect 964 496 994 522
rect 1052 496 1082 522
rect 1140 496 1170 522
rect 1230 496 1260 522
rect 1318 496 1348 522
rect 81 270 111 312
rect 168 270 198 312
rect 256 270 286 312
rect 344 270 374 312
rect 44 251 374 270
rect 44 217 60 251
rect 358 217 374 251
rect 44 204 374 217
rect 81 179 111 204
rect 168 179 198 204
rect 256 179 286 204
rect 344 179 374 204
rect 432 270 462 312
rect 524 270 554 312
rect 612 270 642 312
rect 700 270 730 312
rect 788 270 818 312
rect 876 270 906 312
rect 964 270 994 312
rect 1052 270 1082 312
rect 1140 270 1170 312
rect 1230 270 1260 312
rect 1318 270 1348 312
rect 432 251 1348 270
rect 432 217 456 251
rect 1328 217 1348 251
rect 432 206 1348 217
rect 432 179 462 206
rect 524 179 554 206
rect 612 179 642 206
rect 700 179 730 206
rect 788 179 818 206
rect 876 179 906 206
rect 964 179 994 206
rect 1052 179 1082 206
rect 1140 179 1170 206
rect 1230 179 1260 206
rect 1318 179 1348 206
rect 81 22 111 48
rect 168 22 198 48
rect 256 22 286 48
rect 344 22 374 48
rect 432 22 462 48
rect 524 22 554 48
rect 612 22 642 48
rect 700 22 730 48
rect 788 22 818 48
rect 876 22 906 48
rect 964 22 994 48
rect 1052 22 1082 48
rect 1140 22 1170 48
rect 1230 22 1260 48
rect 1318 22 1348 48
<< polycont >>
rect 60 217 358 251
rect 456 217 1328 251
<< locali >>
rect 0 561 1472 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 526 1472 527
rect 36 480 70 526
rect 36 378 70 394
rect 122 476 156 492
rect 210 482 244 526
rect 210 391 244 407
rect 298 476 332 492
rect 122 357 156 360
rect 386 484 420 526
rect 386 392 420 408
rect 478 476 512 492
rect 298 357 332 360
rect 122 323 444 357
rect 38 251 374 289
rect 38 217 60 251
rect 358 217 374 251
rect 38 214 374 217
rect 410 270 444 323
rect 566 484 600 526
rect 566 393 600 409
rect 654 476 688 492
rect 512 322 654 340
rect 478 320 654 322
rect 742 484 776 526
rect 742 393 776 409
rect 830 476 864 492
rect 688 320 830 340
rect 918 484 952 526
rect 918 393 952 409
rect 1006 476 1040 492
rect 864 320 1006 340
rect 1094 484 1128 526
rect 1094 393 1128 409
rect 1184 476 1218 492
rect 1040 320 1184 340
rect 1272 484 1306 526
rect 1272 393 1306 409
rect 1360 476 1394 492
rect 1218 320 1360 340
rect 1394 320 1444 359
rect 478 306 1444 320
rect 410 251 1344 270
rect 410 217 456 251
rect 1328 217 1344 251
rect 410 180 444 217
rect 1378 183 1444 306
rect 122 150 444 180
rect 36 132 70 148
rect 36 21 70 64
rect 156 146 298 150
rect 122 56 156 72
rect 194 98 260 112
rect 194 64 210 98
rect 244 64 260 98
rect 194 62 260 64
rect 332 146 444 150
rect 478 162 1444 183
rect 478 150 1406 162
rect 210 21 244 62
rect 298 56 332 72
rect 370 98 436 112
rect 370 64 386 98
rect 420 64 436 98
rect 370 62 436 64
rect 512 149 654 150
rect 386 21 420 62
rect 478 56 512 72
rect 566 99 600 115
rect 566 21 600 64
rect 688 149 830 150
rect 654 56 688 72
rect 742 95 776 115
rect 742 21 776 60
rect 864 149 1006 150
rect 830 56 864 72
rect 918 95 952 115
rect 918 21 952 60
rect 1040 149 1182 150
rect 1006 56 1040 72
rect 1094 99 1128 115
rect 1094 21 1128 58
rect 1216 149 1360 150
rect 1182 56 1216 72
rect 1272 99 1306 115
rect 1272 21 1306 58
rect 1394 149 1406 150
rect 1360 56 1394 72
rect 0 17 1472 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_11
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 170 255 204 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 187 272 187 272 0 FreeSans 200 0 0 0 A
flabel locali s 255 255 289 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 272 272 272 272 0 FreeSans 200 0 0 0 A
flabel locali s 68 255 102 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 1394 306 1428 340 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 1411 323 1411 323 0 FreeSans 200 0 0 0 Y
flabel locali s 1394 187 1428 221 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 1411 204 1411 204 0 FreeSans 200 0 0 0 Y
flabel locali s 85 272 85 272 0 FreeSans 200 0 0 0 A
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_11.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1472 220
string MASKHINTS_NSDM 0 -38 1472 204
string MASKHINTS_PSDM 0 287 1472 582
<< end >>
