magic
tech sky130A
magscale 1 2
timestamp 1749429620
<< nwell >>
rect -38 262 1142 582
<< pwell >>
rect 0 28 1104 204
rect 0 26 828 28
rect 22 24 90 26
rect 22 22 110 24
rect 168 22 198 24
rect 256 22 286 24
rect 344 22 374 24
rect 432 22 462 24
rect 519 22 549 24
rect 605 22 635 24
rect 691 22 721 24
rect 784 22 814 24
rect 872 22 902 24
rect 958 22 988 24
rect 22 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 168 298 198 496
rect 256 298 286 496
rect 344 298 374 496
rect 432 298 462 496
rect 519 298 549 496
rect 605 298 635 496
rect 691 298 721 496
rect 784 298 814 496
rect 872 298 902 496
rect 958 298 988 496
<< nmoslvt >>
rect 80 48 110 178
rect 168 48 198 178
rect 256 48 286 178
rect 344 48 374 178
rect 432 48 462 178
rect 519 48 549 178
rect 605 48 635 178
rect 691 48 721 178
rect 784 48 814 178
rect 872 48 902 178
rect 958 48 988 178
<< ndiff >>
rect 27 140 80 178
rect 27 76 35 140
rect 69 76 80 140
rect 27 48 80 76
rect 110 170 168 178
rect 110 72 121 170
rect 155 72 168 170
rect 110 48 168 72
rect 198 170 256 178
rect 198 58 209 170
rect 243 58 256 170
rect 198 48 256 58
rect 286 170 344 178
rect 286 72 298 170
rect 332 72 344 170
rect 286 48 344 72
rect 374 106 432 178
rect 374 72 386 106
rect 420 72 432 106
rect 374 48 432 72
rect 462 170 519 178
rect 462 72 474 170
rect 508 72 519 170
rect 462 48 519 72
rect 549 166 605 178
rect 549 57 560 166
rect 594 57 605 166
rect 549 48 605 57
rect 635 160 691 178
rect 635 126 646 160
rect 680 126 691 160
rect 635 48 691 126
rect 721 170 784 178
rect 721 57 736 170
rect 770 57 784 170
rect 721 48 784 57
rect 814 158 872 178
rect 814 124 826 158
rect 860 124 872 158
rect 814 48 872 124
rect 902 170 958 178
rect 902 58 913 170
rect 947 58 958 170
rect 902 48 958 58
rect 988 156 1077 178
rect 988 122 1002 156
rect 1036 122 1077 156
rect 988 48 1077 122
<< pdiff >>
rect 27 484 80 496
rect 27 350 35 484
rect 69 350 80 484
rect 27 298 80 350
rect 110 476 168 496
rect 110 331 121 476
rect 155 331 168 476
rect 110 298 168 331
rect 198 488 256 496
rect 198 346 209 488
rect 243 346 256 488
rect 198 298 256 346
rect 286 476 344 496
rect 286 354 298 476
rect 332 354 344 476
rect 286 298 344 354
rect 374 474 432 496
rect 374 354 386 474
rect 420 354 432 474
rect 374 298 432 354
rect 462 474 519 496
rect 462 354 474 474
rect 508 354 519 474
rect 462 298 519 354
rect 549 488 605 496
rect 549 342 560 488
rect 594 342 605 488
rect 549 298 605 342
rect 635 474 691 496
rect 635 331 646 474
rect 680 331 691 474
rect 635 298 691 331
rect 721 488 784 496
rect 721 342 734 488
rect 768 342 784 488
rect 721 298 784 342
rect 814 474 872 496
rect 814 331 826 474
rect 860 331 872 474
rect 814 298 872 331
rect 902 488 958 496
rect 902 346 913 488
rect 947 346 958 488
rect 902 298 958 346
rect 988 476 1077 496
rect 988 332 1002 476
rect 1036 332 1077 476
rect 988 298 1077 332
<< ndiffc >>
rect 35 76 69 140
rect 121 72 155 170
rect 209 58 243 170
rect 298 72 332 170
rect 386 72 420 106
rect 474 72 508 170
rect 560 57 594 166
rect 646 126 680 160
rect 736 57 770 170
rect 826 124 860 158
rect 913 58 947 170
rect 1002 122 1036 156
<< pdiffc >>
rect 35 350 69 484
rect 121 331 155 476
rect 209 346 243 488
rect 298 354 332 476
rect 386 354 420 474
rect 474 354 508 474
rect 560 342 594 488
rect 646 331 680 474
rect 734 342 768 488
rect 826 331 860 474
rect 913 346 947 488
rect 1002 332 1036 476
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 519 496 549 522
rect 605 496 635 522
rect 691 496 721 522
rect 784 496 814 522
rect 872 496 902 522
rect 958 496 988 522
rect 80 282 110 298
rect 168 282 198 298
rect 80 268 198 282
rect 256 268 286 298
rect 344 282 374 298
rect 432 282 462 298
rect 519 282 549 298
rect 605 282 635 298
rect 691 282 721 298
rect 784 282 814 298
rect 872 282 902 298
rect 958 282 988 298
rect 344 268 988 282
rect 80 260 286 268
rect 36 250 286 260
rect 36 216 52 250
rect 86 226 286 250
rect 86 216 110 226
rect 36 196 110 216
rect 80 178 110 196
rect 168 178 198 226
rect 256 178 286 226
rect 328 250 988 268
rect 328 216 338 250
rect 372 232 988 250
rect 372 216 390 232
rect 328 200 390 216
rect 344 178 374 200
rect 432 178 462 232
rect 519 178 549 232
rect 605 178 635 232
rect 691 178 721 232
rect 784 178 814 232
rect 872 178 902 232
rect 958 178 988 232
rect 80 22 110 48
rect 168 22 198 48
rect 256 22 286 48
rect 344 22 374 48
rect 432 22 462 48
rect 519 22 549 48
rect 605 22 635 48
rect 691 22 721 48
rect 784 22 814 48
rect 872 22 902 48
rect 958 22 988 48
<< polycont >>
rect 52 216 86 250
rect 338 216 372 250
<< locali >>
rect 0 561 1104 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 526 1104 527
rect 35 484 69 526
rect 35 334 69 350
rect 120 476 156 492
rect 120 331 121 476
rect 155 331 156 476
rect 34 250 86 300
rect 34 216 52 250
rect 34 198 86 216
rect 120 284 156 331
rect 209 488 243 526
rect 209 330 243 346
rect 298 476 332 492
rect 298 284 332 354
rect 386 474 420 526
rect 386 338 420 354
rect 474 474 508 490
rect 474 304 508 354
rect 560 488 594 526
rect 560 326 594 342
rect 646 474 680 490
rect 120 268 332 284
rect 424 292 508 304
rect 646 292 680 331
rect 734 488 768 526
rect 734 326 768 342
rect 826 474 860 490
rect 826 292 860 331
rect 913 488 947 526
rect 913 326 947 346
rect 1002 476 1042 492
rect 1036 332 1042 476
rect 1002 292 1042 332
rect 120 250 378 268
rect 120 244 338 250
rect 120 170 156 244
rect 298 216 338 244
rect 372 216 378 250
rect 424 248 1042 292
rect 424 226 508 248
rect 298 200 378 216
rect 35 140 69 158
rect 35 21 69 76
rect 120 72 121 170
rect 155 72 156 170
rect 120 56 156 72
rect 209 170 243 192
rect 209 21 243 58
rect 298 170 332 200
rect 474 170 508 226
rect 298 56 332 72
rect 386 106 420 122
rect 386 21 420 72
rect 474 56 508 72
rect 560 166 594 182
rect 646 160 680 248
rect 826 244 1042 248
rect 646 110 680 126
rect 736 170 770 190
rect 560 21 594 57
rect 826 158 860 244
rect 826 108 860 124
rect 913 170 947 190
rect 736 21 770 57
rect 1002 156 1042 244
rect 1036 122 1042 156
rect 1002 106 1042 122
rect 913 21 947 58
rect 0 17 1104 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_8
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1104 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali 425 255 459 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 442 272 442 272 0 FreeSans 200 0 0 0 Y
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_8.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1104 216
string MASKHINTS_NSDM 0 -38 1104 204
string MASKHINTS_PSDM 0 272 1104 582
<< end >>
