magic
tech sky130A
magscale 1 2
timestamp 1737034163
<< nwell >>
rect -38 262 314 582
<< pwell >>
rect 0 22 276 204
rect 26 -15 76 22
rect 26 -20 66 -15
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
<< nmoslvt >>
rect 80 49 110 178
rect 166 49 196 178
<< ndiff >>
rect 27 150 80 178
rect 27 62 35 150
rect 69 62 80 150
rect 27 49 80 62
rect 110 170 166 178
rect 110 72 121 170
rect 155 72 166 170
rect 110 49 166 72
rect 196 166 249 178
rect 196 61 207 166
rect 241 61 249 166
rect 196 49 249 61
<< pdiff >>
rect 27 484 80 496
rect 27 318 35 484
rect 69 318 80 484
rect 27 298 80 318
rect 110 476 166 496
rect 110 306 121 476
rect 155 306 166 476
rect 110 298 166 306
rect 196 484 249 496
rect 196 318 207 484
rect 241 318 249 484
rect 196 298 249 318
<< ndiffc >>
rect 35 62 69 150
rect 121 72 155 170
rect 207 61 241 166
<< pdiffc >>
rect 35 318 69 484
rect 121 306 155 476
rect 207 318 241 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 80 268 110 298
rect 166 268 196 298
rect 30 250 196 268
rect 30 216 46 250
rect 80 216 196 250
rect 30 200 196 216
rect 80 178 110 200
rect 166 178 196 200
rect 80 23 110 49
rect 166 23 196 49
<< polycont >>
rect 46 216 80 250
<< locali >>
rect 0 561 276 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 526 276 527
rect 35 484 69 526
rect 35 302 69 318
rect 114 476 158 492
rect 114 306 121 476
rect 155 306 158 476
rect 30 250 80 268
rect 30 216 46 250
rect 30 200 80 216
rect 114 170 158 306
rect 206 484 242 526
rect 206 318 207 484
rect 241 318 242 484
rect 206 302 242 318
rect 35 150 69 166
rect 35 21 69 62
rect 114 72 121 170
rect 155 72 158 170
rect 114 56 158 72
rect 206 166 242 188
rect 206 61 207 166
rect 241 61 242 166
rect 206 21 242 61
rect 0 17 276 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 276 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 276 48 1 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali 34 221 68 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 51 238 51 238 0 FreeSans 200 0 0 0 A
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 276 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__inv_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 276 214
string MASKHINTS_NSDM 0 -38 276 204
string MASKHINTS_PSDM 0 272 276 582
<< end >>
