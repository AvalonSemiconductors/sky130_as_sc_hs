magic
tech sky130A
magscale 1 2
timestamp 1740066495
<< nwell >>
rect -38 262 682 582
<< pwell >>
rect 0 28 644 204
rect 0 22 460 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 338 298 368 496
rect 424 298 454 496
rect 510 298 540 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 252 48 282 178
rect 338 48 368 178
rect 424 48 454 178
rect 510 48 540 178
<< ndiff >>
rect 27 148 80 178
rect 27 72 35 148
rect 69 72 80 148
rect 27 48 80 72
rect 110 90 166 178
rect 110 56 121 90
rect 155 56 166 90
rect 110 48 166 56
rect 196 148 252 178
rect 196 72 207 148
rect 241 72 252 148
rect 196 48 252 72
rect 282 90 338 178
rect 282 56 293 90
rect 327 56 338 90
rect 282 48 338 56
rect 368 148 424 178
rect 368 72 379 148
rect 413 72 424 148
rect 368 48 424 72
rect 454 162 510 178
rect 454 128 465 162
rect 499 128 510 162
rect 454 48 510 128
rect 540 90 617 178
rect 540 56 551 90
rect 585 56 617 90
rect 540 48 617 56
<< pdiff >>
rect 27 484 80 496
rect 27 398 35 484
rect 69 398 80 484
rect 27 298 80 398
rect 110 488 166 496
rect 110 454 121 488
rect 155 454 166 488
rect 110 298 166 454
rect 196 402 252 496
rect 196 368 207 402
rect 241 368 252 402
rect 196 298 252 368
rect 282 488 338 496
rect 282 454 293 488
rect 327 454 338 488
rect 282 298 338 454
rect 368 486 424 496
rect 368 452 379 486
rect 413 452 424 486
rect 368 298 424 452
rect 454 476 510 496
rect 454 392 465 476
rect 499 392 510 476
rect 454 298 510 392
rect 540 486 617 496
rect 540 452 551 486
rect 585 452 617 486
rect 540 298 617 452
<< ndiffc >>
rect 35 72 69 148
rect 121 56 155 90
rect 207 72 241 148
rect 293 56 327 90
rect 379 72 413 148
rect 465 128 499 162
rect 551 56 585 90
<< pdiffc >>
rect 35 398 69 484
rect 121 454 155 488
rect 207 368 241 402
rect 293 454 327 488
rect 379 452 413 486
rect 465 392 499 476
rect 551 452 585 486
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 424 496 454 522
rect 510 496 540 522
rect 80 270 110 298
rect 44 250 110 270
rect 44 216 58 250
rect 92 216 110 250
rect 44 198 110 216
rect 80 178 110 198
rect 166 270 196 298
rect 252 270 282 298
rect 338 270 368 298
rect 424 270 454 298
rect 510 270 540 298
rect 166 250 282 270
rect 166 216 202 250
rect 236 216 282 250
rect 166 198 282 216
rect 324 250 378 270
rect 324 216 334 250
rect 368 216 378 250
rect 324 198 378 216
rect 420 250 540 270
rect 420 216 430 250
rect 464 216 540 250
rect 420 198 540 216
rect 166 178 196 198
rect 252 178 282 198
rect 338 178 368 198
rect 424 178 454 198
rect 510 178 540 198
rect 80 22 110 48
rect 166 22 196 48
rect 252 22 282 48
rect 338 22 368 48
rect 424 22 454 48
rect 510 22 540 48
<< polycont >>
rect 58 216 92 250
rect 202 216 236 250
rect 334 216 368 250
rect 430 216 464 250
<< locali >>
rect 0 561 644 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 526 644 527
rect 35 484 69 526
rect 104 454 121 488
rect 155 454 293 488
rect 327 454 345 488
rect 379 486 413 526
rect 379 436 413 452
rect 465 476 499 492
rect 35 376 69 398
rect 191 368 207 402
rect 241 392 465 402
rect 551 486 585 526
rect 551 436 585 452
rect 499 392 542 402
rect 241 368 542 392
rect 508 348 542 368
rect 44 300 372 334
rect 44 250 94 300
rect 324 270 372 300
rect 420 270 466 334
rect 44 216 58 250
rect 92 216 94 250
rect 44 198 94 216
rect 166 250 282 266
rect 166 216 202 250
rect 236 216 282 250
rect 166 202 282 216
rect 324 250 378 270
rect 324 216 334 250
rect 368 216 378 250
rect 324 198 378 216
rect 420 250 474 270
rect 420 216 430 250
rect 464 216 474 250
rect 420 198 474 216
rect 508 200 566 348
rect 35 148 413 164
rect 508 162 542 200
rect 69 130 207 148
rect 35 56 69 72
rect 104 56 121 90
rect 155 56 172 90
rect 241 130 379 148
rect 207 56 241 72
rect 276 56 293 90
rect 327 56 344 90
rect 448 128 465 162
rect 499 128 542 162
rect 413 72 551 90
rect 379 56 551 72
rect 585 56 602 90
rect 121 21 155 56
rect 293 21 327 56
rect 0 17 644 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel comment s 0 0 0 0 4 oai21_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 51 204 85 238 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 68 221 68 221 0 FreeSans 200 0 0 0 A
flabel locali s 221 204 255 238 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 238 221 238 221 0 FreeSans 200 0 0 0 B
flabel locali s 425 204 459 238 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 442 221 442 221 0 FreeSans 200 0 0 0 C
flabel locali s 527 204 561 238 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 544 221 544 221 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__oai21_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 644 220
string MASKHINTS_NSDM 0 -38 644 209
string MASKHINTS_PSDM 0 273 644 582
<< end >>
