magic
tech sky130A
magscale 1 2
timestamp 1738754271
<< nwell >>
rect -38 262 958 582
<< pwell >>
rect 0 24 920 204
rect 0 22 736 24
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 338 298 368 496
rect 528 298 558 496
rect 614 298 644 496
rect 700 298 730 496
rect 786 298 816 496
<< nmoslvt >>
rect 80 49 110 178
rect 166 49 196 178
rect 252 49 282 178
rect 338 49 368 178
rect 528 49 558 178
rect 614 49 644 178
rect 700 49 730 178
rect 786 49 816 178
<< ndiff >>
rect 27 106 80 178
rect 27 72 35 106
rect 69 72 80 106
rect 27 49 80 72
rect 110 92 166 178
rect 110 58 121 92
rect 155 58 166 92
rect 110 49 166 58
rect 196 106 252 178
rect 196 72 207 106
rect 241 72 252 106
rect 196 49 252 72
rect 282 170 338 178
rect 282 136 293 170
rect 327 136 338 170
rect 282 49 338 136
rect 368 106 421 178
rect 368 72 379 106
rect 413 72 421 106
rect 368 49 421 72
rect 475 96 528 178
rect 475 62 483 96
rect 517 62 528 96
rect 475 49 528 62
rect 558 170 614 178
rect 558 71 569 170
rect 603 71 614 170
rect 558 49 614 71
rect 644 94 700 178
rect 644 60 655 94
rect 689 60 700 94
rect 644 49 700 60
rect 730 164 786 178
rect 730 72 741 164
rect 775 72 786 164
rect 730 49 786 72
rect 816 166 873 178
rect 816 57 827 166
rect 861 57 873 166
rect 816 49 873 57
<< pdiff >>
rect 27 476 80 496
rect 27 348 35 476
rect 69 348 80 476
rect 27 298 80 348
rect 110 476 166 496
rect 110 340 121 476
rect 155 340 166 476
rect 110 298 166 340
rect 196 488 252 496
rect 196 408 207 488
rect 241 408 252 488
rect 196 298 252 408
rect 282 476 338 496
rect 282 324 293 476
rect 327 324 338 476
rect 282 298 338 324
rect 368 484 421 496
rect 368 408 379 484
rect 413 408 421 484
rect 368 298 421 408
rect 475 474 528 496
rect 475 408 483 474
rect 517 408 528 474
rect 475 298 528 408
rect 558 406 614 496
rect 558 324 569 406
rect 603 324 614 406
rect 558 298 614 324
rect 644 488 700 496
rect 644 384 655 488
rect 689 384 700 488
rect 644 298 700 384
rect 730 406 786 496
rect 730 316 741 406
rect 775 316 786 406
rect 730 298 786 316
rect 816 474 869 496
rect 816 342 827 474
rect 861 342 869 474
rect 816 298 869 342
<< ndiffc >>
rect 35 72 69 106
rect 121 58 155 92
rect 207 72 241 106
rect 293 136 327 170
rect 379 72 413 106
rect 483 62 517 96
rect 569 71 603 170
rect 655 60 689 94
rect 741 72 775 164
rect 827 57 861 166
<< pdiffc >>
rect 35 348 69 476
rect 121 340 155 476
rect 207 408 241 488
rect 293 324 327 476
rect 379 408 413 484
rect 483 408 517 474
rect 569 324 603 406
rect 655 384 689 488
rect 741 316 775 406
rect 827 342 861 474
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 528 496 558 522
rect 614 496 644 522
rect 700 496 730 522
rect 786 496 816 522
rect 80 274 110 298
rect 166 274 196 298
rect 64 250 196 274
rect 64 216 80 250
rect 114 216 196 250
rect 64 206 196 216
rect 80 178 110 206
rect 166 178 196 206
rect 252 276 282 298
rect 338 276 368 298
rect 252 250 368 276
rect 252 216 268 250
rect 302 216 368 250
rect 252 206 368 216
rect 252 178 282 206
rect 338 178 368 206
rect 528 276 558 298
rect 614 276 644 298
rect 528 250 644 276
rect 528 216 544 250
rect 578 216 644 250
rect 528 206 644 216
rect 528 178 558 206
rect 614 178 644 206
rect 700 276 730 298
rect 786 276 816 298
rect 700 250 846 276
rect 700 216 796 250
rect 830 216 846 250
rect 700 206 846 216
rect 700 178 730 206
rect 786 178 816 206
rect 80 23 110 49
rect 166 23 196 49
rect 252 23 282 49
rect 338 23 368 49
rect 528 23 558 49
rect 614 23 644 49
rect 700 23 730 49
rect 786 23 816 49
<< polycont >>
rect 80 216 114 250
rect 268 216 302 250
rect 544 216 578 250
rect 796 216 830 250
<< locali >>
rect 0 561 920 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 526 920 527
rect 30 476 74 526
rect 30 348 35 476
rect 69 348 74 476
rect 30 332 74 348
rect 118 476 158 492
rect 118 340 121 476
rect 155 358 158 476
rect 202 488 246 526
rect 202 408 207 488
rect 241 408 246 488
rect 202 392 246 408
rect 290 476 330 492
rect 290 358 293 476
rect 155 340 293 358
rect 118 324 293 340
rect 327 358 330 476
rect 374 484 418 526
rect 374 408 379 484
rect 413 408 418 484
rect 374 392 418 408
rect 480 488 864 490
rect 480 474 655 488
rect 480 408 483 474
rect 517 456 655 474
rect 517 408 520 456
rect 480 392 520 408
rect 566 406 608 422
rect 566 358 569 406
rect 327 324 569 358
rect 603 324 608 406
rect 650 384 655 456
rect 689 474 864 488
rect 689 456 827 474
rect 689 384 694 456
rect 650 368 694 384
rect 740 406 780 422
rect 740 334 741 406
rect 118 322 608 324
rect 566 308 608 322
rect 692 316 741 334
rect 775 316 780 406
rect 824 342 827 456
rect 861 342 864 474
rect 824 326 864 342
rect 692 300 780 316
rect 64 250 196 266
rect 64 216 80 250
rect 114 216 196 250
rect 252 250 390 266
rect 252 216 268 250
rect 302 216 390 250
rect 492 250 644 266
rect 492 216 544 250
rect 578 216 644 250
rect 692 182 746 300
rect 780 250 858 266
rect 780 216 796 250
rect 830 216 858 250
rect 32 142 242 178
rect 32 106 74 142
rect 32 72 35 106
rect 69 72 74 106
rect 32 56 74 72
rect 116 92 160 108
rect 116 58 121 92
rect 155 58 160 92
rect 116 21 160 58
rect 202 106 242 142
rect 276 170 786 182
rect 276 136 293 170
rect 327 146 569 170
rect 327 136 344 146
rect 202 72 207 106
rect 241 96 242 106
rect 362 96 379 106
rect 241 72 379 96
rect 413 72 430 106
rect 202 56 430 72
rect 478 96 522 112
rect 478 62 483 96
rect 517 62 522 96
rect 478 21 522 62
rect 566 71 569 146
rect 603 164 786 170
rect 603 146 741 164
rect 603 71 606 146
rect 566 56 606 71
rect 650 94 694 112
rect 650 60 655 94
rect 689 60 694 94
rect 569 55 603 56
rect 650 21 694 60
rect 738 72 741 146
rect 775 72 786 164
rect 738 55 786 72
rect 824 166 864 182
rect 824 57 827 166
rect 861 57 864 166
rect 824 21 864 57
rect 0 17 920 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 aoi211_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 85 221 119 255 0 FreeSans 200 0 0 0 A
port 9 nsew signal input
flabel locali 102 238 102 238 0 FreeSans 200 0 0 0 A
flabel locali 272 221 306 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 289 238 289 238 0 FreeSans 200 0 0 0 B
flabel locali 544 221 578 255 0 FreeSans 200 0 0 0 C
port 6 nsew signal input
flabel locali 561 238 561 238 0 FreeSans 200 0 0 0 C
flabel locali 799 221 833 255 0 FreeSans 200 0 0 1 D
port 7 nsew signal input
flabel locali 816 238 816 238 0 FreeSans 200 0 0 1 D
flabel locali 697 221 731 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali 714 238 714 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__aoi211_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 920 214
string MASKHINTS_NSDM 0 -38 920 204
string MASKHINTS_PSDM 0 272 920 582
<< end >>
