magic
tech sky130A
magscale 1 2
timestamp 1740057465
<< nwell >>
rect -38 262 866 582
<< pwell >>
rect 0 28 828 204
rect 0 22 736 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 404 298 434 496
rect 602 298 632 496
rect 688 298 718 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 252 48 282 178
rect 404 48 434 178
rect 602 48 632 178
rect 688 48 718 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 92 166 178
rect 110 58 121 92
rect 155 58 166 92
rect 110 48 166 58
rect 196 150 252 178
rect 196 72 207 150
rect 241 72 252 150
rect 196 48 252 72
rect 282 166 404 178
rect 282 132 302 166
rect 336 132 404 166
rect 282 48 404 132
rect 434 90 491 178
rect 434 56 445 90
rect 479 56 491 90
rect 434 48 491 56
rect 545 92 602 178
rect 545 58 557 92
rect 591 58 602 92
rect 545 48 602 58
rect 632 170 688 178
rect 632 72 643 170
rect 677 72 688 170
rect 632 48 688 72
rect 718 150 801 178
rect 718 56 729 150
rect 763 56 801 150
rect 718 48 801 56
<< pdiff >>
rect 27 480 80 496
rect 27 444 35 480
rect 69 444 80 480
rect 27 298 80 444
rect 110 298 166 496
rect 196 476 252 496
rect 196 426 207 476
rect 241 426 252 476
rect 196 298 252 426
rect 282 298 404 496
rect 434 488 602 496
rect 434 334 446 488
rect 591 334 602 488
rect 434 298 602 334
rect 632 476 688 496
rect 632 306 643 476
rect 677 306 688 476
rect 632 298 688 306
rect 718 488 801 496
rect 718 338 729 488
rect 763 338 801 488
rect 718 298 801 338
<< ndiffc >>
rect 35 72 69 150
rect 121 58 155 92
rect 207 72 241 150
rect 302 132 336 166
rect 445 56 479 90
rect 557 58 591 92
rect 643 72 677 170
rect 729 56 763 150
<< pdiffc >>
rect 35 444 69 480
rect 207 426 241 476
rect 446 334 591 488
rect 643 306 677 476
rect 729 338 763 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 404 496 434 522
rect 602 496 632 522
rect 688 496 718 522
rect 80 266 110 298
rect 166 266 196 298
rect 252 266 282 298
rect 404 266 434 298
rect 602 268 632 298
rect 688 268 718 298
rect 56 250 110 266
rect 56 216 66 250
rect 100 216 110 250
rect 56 200 110 216
rect 152 250 206 266
rect 152 216 162 250
rect 196 216 206 250
rect 152 200 206 216
rect 248 250 302 266
rect 248 216 258 250
rect 292 216 302 250
rect 248 200 302 216
rect 404 250 458 266
rect 404 216 414 250
rect 448 216 458 250
rect 80 178 110 200
rect 166 178 196 200
rect 252 178 282 200
rect 404 198 458 216
rect 554 250 718 268
rect 554 216 564 250
rect 598 216 718 250
rect 554 200 718 216
rect 404 178 434 198
rect 602 178 632 200
rect 688 178 718 200
rect 80 22 110 48
rect 166 22 196 48
rect 252 22 282 48
rect 404 22 434 48
rect 602 22 632 48
rect 688 22 718 48
<< polycont >>
rect 66 216 100 250
rect 162 216 196 250
rect 258 216 292 250
rect 414 216 448 250
rect 564 216 598 250
<< locali >>
rect 0 561 828 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 526 828 527
rect 35 480 69 526
rect 35 428 69 444
rect 207 476 241 492
rect 446 488 592 526
rect 241 426 370 444
rect 207 410 370 426
rect 38 266 88 394
rect 144 266 186 382
rect 240 266 290 376
rect 38 250 110 266
rect 38 216 66 250
rect 100 216 110 250
rect 38 200 110 216
rect 144 250 206 266
rect 144 216 162 250
rect 196 216 206 250
rect 144 200 206 216
rect 240 250 302 266
rect 240 216 258 250
rect 292 216 302 250
rect 240 200 302 216
rect 35 150 241 166
rect 69 132 207 150
rect 35 56 69 72
rect 104 58 121 92
rect 155 58 172 92
rect 286 132 302 166
rect 336 160 370 410
rect 591 334 592 488
rect 446 318 592 334
rect 643 476 677 492
rect 729 488 763 526
rect 729 322 763 338
rect 643 294 677 306
rect 404 250 490 284
rect 404 216 414 250
rect 448 216 490 250
rect 404 194 490 216
rect 544 250 608 268
rect 544 216 564 250
rect 598 216 608 250
rect 544 200 608 216
rect 544 160 578 200
rect 336 132 578 160
rect 286 126 578 132
rect 643 194 708 294
rect 643 170 677 194
rect 241 72 445 90
rect 121 21 155 58
rect 207 56 445 72
rect 479 56 495 90
rect 540 58 557 92
rect 591 58 608 92
rect 557 21 591 58
rect 643 56 677 72
rect 729 150 763 166
rect 729 21 763 56
rect 0 17 828 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel comment s 0 0 0 0 4 oa22_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 68 221 102 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 85 238 85 238 0 FreeSans 200 0 0 0 A
flabel locali s 153 221 187 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 170 238 170 238 0 FreeSans 200 0 0 0 B
flabel locali s 255 221 289 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 272 238 272 238 0 FreeSans 200 0 0 0 C
flabel locali s 442 221 476 255 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel locali s 459 238 459 238 0 FreeSans 200 0 0 0 D
flabel locali s 663 221 697 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 680 238 680 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__oa22_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 828 220
string MASKHINTS_NSDM 0 -38 828 209
string MASKHINTS_PSDM 0 273 828 582
<< end >>
