magic
tech sky130A
magscale 1 2
timestamp 1738771478
<< nwell >>
rect -38 262 1786 582
<< pwell >>
rect 18 48 1742 204
rect 22 44 1608 48
rect 22 -15 82 44
rect 22 -20 64 -15
<< pmos >>
rect 83 331 113 496
rect 170 331 200 496
rect 368 388 398 496
rect 466 412 496 496
rect 584 412 614 496
rect 754 402 784 496
rect 854 402 884 496
rect 962 410 992 496
rect 1080 410 1110 496
rect 1250 402 1280 496
rect 1352 402 1382 496
rect 1542 298 1572 496
rect 1628 298 1658 496
<< nmoslvt >>
rect 83 49 113 162
rect 170 49 200 162
rect 368 49 398 164
rect 468 49 498 138
rect 582 49 612 138
rect 754 49 784 138
rect 854 49 884 148
rect 964 49 994 144
rect 1076 49 1106 144
rect 1250 49 1280 144
rect 1352 49 1382 144
rect 1542 49 1572 178
rect 1628 49 1658 178
<< ndiff >>
rect 30 128 83 162
rect 30 72 38 128
rect 72 72 83 128
rect 30 49 83 72
rect 113 112 170 162
rect 113 60 124 112
rect 158 60 170 112
rect 113 49 170 60
rect 200 134 258 162
rect 200 72 212 134
rect 246 72 258 134
rect 200 49 258 72
rect 312 122 368 164
rect 312 64 322 122
rect 356 64 368 122
rect 312 49 368 64
rect 398 138 448 164
rect 804 138 854 148
rect 398 130 468 138
rect 398 72 416 130
rect 450 72 468 130
rect 398 49 468 72
rect 498 120 582 138
rect 498 86 526 120
rect 560 86 582 120
rect 498 49 582 86
rect 612 49 754 138
rect 784 114 854 138
rect 784 60 806 114
rect 840 60 854 114
rect 784 49 854 60
rect 884 144 942 148
rect 1489 150 1542 178
rect 884 130 964 144
rect 884 74 910 130
rect 944 74 964 130
rect 884 49 964 74
rect 994 120 1076 144
rect 994 86 1022 120
rect 1056 86 1076 120
rect 994 49 1076 86
rect 1106 49 1250 144
rect 1280 114 1352 144
rect 1280 60 1304 114
rect 1338 60 1352 114
rect 1280 49 1352 60
rect 1382 138 1434 144
rect 1382 126 1435 138
rect 1382 72 1393 126
rect 1427 72 1435 126
rect 1382 49 1435 72
rect 1489 68 1497 150
rect 1531 68 1542 150
rect 1489 49 1542 68
rect 1572 158 1628 178
rect 1572 80 1583 158
rect 1617 80 1628 158
rect 1572 49 1628 80
rect 1658 166 1711 178
rect 1658 68 1669 166
rect 1703 68 1711 166
rect 1658 49 1711 68
<< pdiff >>
rect 28 470 83 496
rect 28 378 38 470
rect 72 378 83 470
rect 28 331 83 378
rect 113 484 170 496
rect 113 434 124 484
rect 158 434 170 484
rect 113 331 170 434
rect 200 470 258 496
rect 200 374 212 470
rect 246 374 258 470
rect 312 484 368 496
rect 312 432 322 484
rect 356 432 368 484
rect 312 388 368 432
rect 398 472 466 496
rect 398 432 416 472
rect 450 432 466 472
rect 398 412 466 432
rect 496 476 584 496
rect 496 442 526 476
rect 560 442 584 476
rect 496 412 584 442
rect 614 412 754 496
rect 398 388 448 412
rect 200 331 258 374
rect 630 402 754 412
rect 784 488 854 496
rect 784 432 798 488
rect 832 432 854 488
rect 784 402 854 432
rect 884 474 962 496
rect 884 420 910 474
rect 944 420 962 474
rect 884 410 962 420
rect 992 476 1080 496
rect 992 442 1022 476
rect 1056 442 1080 476
rect 992 410 1080 442
rect 1110 410 1250 496
rect 884 402 934 410
rect 1126 402 1250 410
rect 1280 488 1352 496
rect 1280 432 1302 488
rect 1336 432 1352 488
rect 1280 402 1352 432
rect 1382 476 1435 496
rect 1382 422 1393 476
rect 1427 422 1435 476
rect 1382 402 1435 422
rect 1489 478 1542 496
rect 1489 388 1497 478
rect 1531 388 1542 478
rect 1489 298 1542 388
rect 1572 468 1628 496
rect 1572 402 1583 468
rect 1617 402 1628 468
rect 1572 298 1628 402
rect 1658 480 1711 496
rect 1658 310 1669 480
rect 1703 310 1711 480
rect 1658 298 1711 310
<< ndiffc >>
rect 38 72 72 128
rect 124 60 158 112
rect 212 72 246 134
rect 322 64 356 122
rect 416 72 450 130
rect 526 86 560 120
rect 806 60 840 114
rect 910 74 944 130
rect 1022 86 1056 120
rect 1304 60 1338 114
rect 1393 72 1427 126
rect 1497 68 1531 150
rect 1583 80 1617 158
rect 1669 68 1703 166
<< pdiffc >>
rect 38 378 72 470
rect 124 434 158 484
rect 212 374 246 470
rect 322 432 356 484
rect 416 432 450 472
rect 526 442 560 476
rect 798 432 832 488
rect 910 420 944 474
rect 1022 442 1056 476
rect 1302 432 1336 488
rect 1393 422 1427 476
rect 1497 388 1531 478
rect 1583 402 1617 468
rect 1669 310 1703 480
<< poly >>
rect 83 496 113 522
rect 170 496 200 522
rect 368 496 398 522
rect 466 496 496 522
rect 584 496 614 522
rect 754 496 784 522
rect 854 496 884 522
rect 962 496 992 522
rect 1080 496 1110 522
rect 1250 496 1280 522
rect 1352 496 1382 522
rect 1542 496 1572 522
rect 1628 496 1658 522
rect 83 300 113 331
rect 32 284 113 300
rect 32 250 42 284
rect 76 250 113 284
rect 32 230 113 250
rect 83 162 113 230
rect 170 296 200 331
rect 368 300 398 388
rect 466 372 496 412
rect 466 362 542 372
rect 466 328 488 362
rect 526 328 542 362
rect 466 318 542 328
rect 170 280 228 296
rect 170 246 180 280
rect 214 246 228 280
rect 316 290 398 300
rect 316 256 332 290
rect 366 256 398 290
rect 584 276 614 412
rect 316 246 398 256
rect 170 230 228 246
rect 170 162 200 230
rect 368 164 398 246
rect 468 260 614 276
rect 468 226 488 260
rect 526 246 614 260
rect 754 262 784 402
rect 854 370 884 402
rect 826 354 884 370
rect 826 320 836 354
rect 874 320 884 354
rect 826 304 884 320
rect 962 372 992 410
rect 962 362 1038 372
rect 962 328 980 362
rect 1018 328 1038 362
rect 962 318 1038 328
rect 754 246 812 262
rect 526 226 542 246
rect 468 216 542 226
rect 654 216 712 232
rect 468 138 498 216
rect 654 196 664 216
rect 582 182 664 196
rect 702 182 712 216
rect 582 166 712 182
rect 754 212 764 246
rect 802 212 812 246
rect 754 196 812 212
rect 582 138 612 166
rect 754 138 784 196
rect 854 148 884 304
rect 1080 276 1110 410
rect 964 260 1110 276
rect 964 226 984 260
rect 1022 246 1110 260
rect 1250 262 1280 402
rect 1352 370 1382 402
rect 1322 354 1382 370
rect 1322 320 1336 354
rect 1372 320 1382 354
rect 1322 304 1382 320
rect 1352 270 1382 304
rect 1542 270 1572 298
rect 1628 270 1658 298
rect 1250 246 1308 262
rect 1022 226 1038 246
rect 964 216 1038 226
rect 1150 216 1208 232
rect 964 144 994 216
rect 1150 196 1160 216
rect 1076 182 1160 196
rect 1198 182 1208 216
rect 1076 166 1208 182
rect 1250 212 1260 246
rect 1298 212 1308 246
rect 1250 196 1308 212
rect 1352 206 1658 270
rect 1352 200 1572 206
rect 1076 144 1106 166
rect 1250 144 1280 196
rect 1352 144 1382 200
rect 1542 178 1572 200
rect 1628 178 1658 206
rect 83 23 113 49
rect 170 23 200 49
rect 368 23 398 49
rect 468 23 498 49
rect 582 23 612 49
rect 754 23 784 49
rect 854 23 884 49
rect 964 23 994 49
rect 1076 23 1106 49
rect 1250 23 1280 49
rect 1352 23 1382 49
rect 1542 23 1572 49
rect 1628 23 1658 49
<< polycont >>
rect 42 250 76 284
rect 488 328 526 362
rect 180 246 214 280
rect 332 256 366 290
rect 488 226 526 260
rect 836 320 874 354
rect 980 328 1018 362
rect 664 182 702 216
rect 764 212 802 246
rect 984 226 1022 260
rect 1336 320 1372 354
rect 1160 182 1198 216
rect 1260 212 1298 246
<< locali >>
rect 0 561 1748 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 526 1748 527
rect 38 470 72 488
rect 124 484 158 526
rect 124 418 158 434
rect 212 470 246 488
rect 72 378 156 384
rect 38 350 156 378
rect 322 484 356 526
rect 322 414 356 432
rect 416 472 450 490
rect 798 488 832 526
rect 510 442 526 476
rect 246 374 282 384
rect 212 360 282 374
rect 212 350 248 360
rect 24 284 88 316
rect 24 250 42 284
rect 76 250 88 284
rect 24 234 88 250
rect 122 296 156 350
rect 242 326 248 350
rect 242 318 282 326
rect 122 280 214 296
rect 122 246 180 280
rect 122 230 214 246
rect 122 196 156 230
rect 248 196 282 318
rect 38 162 156 196
rect 212 162 282 196
rect 316 290 382 336
rect 316 256 332 290
rect 366 256 382 290
rect 316 184 382 256
rect 38 128 72 162
rect 212 134 246 162
rect 38 56 72 72
rect 124 112 158 128
rect 124 21 158 60
rect 212 56 246 72
rect 322 122 356 150
rect 322 21 356 64
rect 416 130 450 432
rect 484 362 526 378
rect 484 328 488 362
rect 484 312 526 328
rect 560 356 594 476
rect 798 416 832 432
rect 910 474 944 490
rect 1302 488 1336 526
rect 1006 442 1022 476
rect 834 356 876 370
rect 560 354 876 356
rect 560 322 836 354
rect 484 260 526 276
rect 484 226 488 260
rect 484 210 526 226
rect 560 176 594 322
rect 834 320 836 322
rect 874 320 876 354
rect 834 304 876 320
rect 760 246 802 262
rect 910 246 944 420
rect 978 362 1020 378
rect 978 328 980 362
rect 1018 328 1020 362
rect 978 312 1020 328
rect 1056 358 1090 476
rect 1302 416 1336 432
rect 1388 476 1440 492
rect 1388 422 1393 476
rect 1427 422 1440 476
rect 1388 406 1440 422
rect 1334 358 1372 370
rect 1056 354 1372 358
rect 1056 324 1336 354
rect 542 142 594 176
rect 660 216 702 232
rect 660 180 664 216
rect 760 212 764 246
rect 802 212 944 246
rect 760 196 802 212
rect 660 166 702 180
rect 542 120 576 142
rect 910 130 944 212
rect 980 260 1022 276
rect 980 226 984 260
rect 980 210 1022 226
rect 1056 176 1090 324
rect 1334 320 1336 324
rect 1334 304 1372 320
rect 1256 246 1298 262
rect 1406 246 1440 406
rect 1497 478 1531 526
rect 1497 372 1531 388
rect 1578 468 1622 484
rect 1578 402 1583 468
rect 1617 402 1622 468
rect 1578 338 1622 402
rect 510 86 526 120
rect 560 86 576 120
rect 806 114 840 130
rect 416 56 450 72
rect 806 21 840 60
rect 1038 142 1090 176
rect 1158 216 1200 232
rect 1158 182 1160 216
rect 1198 182 1200 216
rect 1256 212 1260 246
rect 1298 212 1440 246
rect 1538 230 1622 338
rect 1669 480 1703 526
rect 1669 294 1703 310
rect 1256 196 1298 212
rect 1158 166 1200 182
rect 1406 158 1440 212
rect 1038 120 1072 142
rect 1391 134 1440 158
rect 1497 150 1531 166
rect 1006 86 1022 120
rect 1056 86 1072 120
rect 1304 114 1338 130
rect 910 58 944 74
rect 1304 21 1338 60
rect 1391 126 1432 134
rect 1391 72 1393 126
rect 1427 72 1432 126
rect 1391 56 1432 72
rect 1497 21 1531 68
rect 1578 158 1622 230
rect 1578 80 1583 158
rect 1617 80 1622 158
rect 1578 60 1622 80
rect 1669 166 1703 182
rect 1669 21 1703 68
rect 0 17 1748 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 248 326 282 360
rect 180 246 214 280
rect 488 328 526 362
rect 488 226 526 260
rect 980 328 1018 362
rect 664 182 702 216
rect 664 180 702 182
rect 984 226 1022 260
rect 1160 182 1198 216
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 234 362 878 368
rect 234 360 488 362
rect 234 326 248 360
rect 282 328 488 360
rect 526 328 878 362
rect 282 326 878 328
rect 234 322 878 326
rect 968 362 1198 368
rect 968 328 980 362
rect 1018 328 1198 362
rect 968 322 1198 328
rect 234 318 294 322
rect 152 280 228 288
rect 152 246 180 280
rect 214 246 228 280
rect 152 238 228 246
rect 476 260 538 268
rect 152 126 180 238
rect 476 226 488 260
rect 526 226 538 260
rect 660 238 704 322
rect 842 264 878 322
rect 994 266 1022 268
rect 972 264 1034 266
rect 842 260 1034 264
rect 476 220 538 226
rect 500 218 538 220
rect 500 128 528 218
rect 658 216 708 238
rect 842 230 984 260
rect 972 226 984 230
rect 1022 226 1034 260
rect 1154 238 1198 322
rect 972 218 1034 226
rect 658 180 664 216
rect 702 180 708 216
rect 994 210 1022 218
rect 1152 216 1206 238
rect 658 164 708 180
rect 1152 182 1160 216
rect 1198 182 1206 216
rect 1152 164 1206 182
rect 1172 128 1200 164
rect 494 126 1200 128
rect 152 98 1200 126
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxfp_2
flabel locali s 29 272 63 306 0 FreeSans 400 0 0 0 CLK
port 5 nsew clock input
flabel locali s 46 289 46 289 0 FreeSans 400 0 0 0 CLK
flabel locali s 329 238 363 272 0 FreeSans 200 0 0 0 D
port 7 nsew signal input
flabel locali s 346 255 346 255 0 FreeSans 200 0 0 0 D
flabel locali s 1569 272 1603 306 0 FreeSans 200 0 0 0 QN
port 6 nsew signal output
flabel locali s 1586 289 1586 289 0 FreeSans 200 0 0 0 QN
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel metal1 s 0 -48 1748 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__dfxfp_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1748 214
string MASKHINTS_NSDM 0 -38 1748 204
string MASKHINTS_PSDM 0 272 1748 582
<< end >>
