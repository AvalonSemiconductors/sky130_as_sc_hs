magic
tech sky130A
magscale 1 2
timestamp 1740314537
<< nwell >>
rect -38 262 406 582
<< pwell >>
rect 6 42 362 204
rect 22 30 90 42
rect 22 22 110 30
rect 22 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 168 298 198 496
rect 256 298 286 496
<< nmoslvt >>
rect 80 48 110 178
rect 168 48 198 178
rect 256 48 286 178
<< ndiff >>
rect 27 140 80 178
rect 27 106 35 140
rect 69 106 80 140
rect 27 48 80 106
rect 110 92 168 178
rect 110 58 121 92
rect 155 58 168 92
rect 110 48 168 58
rect 198 122 256 178
rect 198 88 210 122
rect 244 88 256 122
rect 198 48 256 88
rect 286 166 340 178
rect 286 64 298 166
rect 332 64 340 166
rect 286 48 340 64
<< pdiff >>
rect 27 466 80 496
rect 27 358 35 466
rect 69 358 80 466
rect 27 298 80 358
rect 110 488 168 496
rect 110 426 121 488
rect 155 426 168 488
rect 110 298 168 426
rect 198 446 256 496
rect 198 412 210 446
rect 244 412 256 446
rect 198 298 256 412
rect 286 482 340 496
rect 286 342 298 482
rect 332 342 340 482
rect 286 298 340 342
<< ndiffc >>
rect 35 106 69 140
rect 121 58 155 92
rect 210 88 244 122
rect 298 64 332 166
<< pdiffc >>
rect 35 358 69 466
rect 121 426 155 488
rect 210 412 244 446
rect 298 342 332 482
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 80 270 110 298
rect 168 272 198 298
rect 50 250 110 270
rect 50 216 66 250
rect 100 216 110 250
rect 50 200 110 216
rect 152 254 206 272
rect 256 254 286 298
rect 152 250 286 254
rect 152 216 162 250
rect 196 224 286 250
rect 196 216 206 224
rect 152 200 206 216
rect 80 178 110 200
rect 168 178 198 200
rect 256 178 286 224
rect 80 22 110 48
rect 168 22 198 48
rect 256 22 286 48
<< polycont >>
rect 66 216 100 250
rect 162 216 196 250
<< locali >>
rect 0 561 368 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 526 368 527
rect 121 488 155 526
rect 35 466 69 484
rect 298 482 332 526
rect 121 410 155 426
rect 210 446 264 462
rect 244 412 264 446
rect 210 396 264 412
rect 69 358 168 376
rect 35 342 168 358
rect 34 250 100 296
rect 34 216 66 250
rect 34 200 100 216
rect 134 274 168 342
rect 230 298 264 396
rect 298 326 332 342
rect 134 250 196 274
rect 134 216 162 250
rect 134 200 196 216
rect 230 246 278 298
rect 134 166 168 200
rect 35 140 168 166
rect 69 132 168 140
rect 230 138 264 246
rect 35 90 69 106
rect 210 122 264 138
rect 104 92 172 98
rect 104 58 121 92
rect 155 58 172 92
rect 244 88 264 122
rect 210 72 264 88
rect 298 166 332 188
rect 121 21 155 58
rect 298 21 332 64
rect 0 17 368 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali s 238 255 272 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 255 272 255 272 0 FreeSans 200 0 0 0 Y
flabel locali s 221 102 255 136 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 238 119 238 119 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 368 216
string MASKHINTS_NSDM 0 -38 368 204
string MASKHINTS_PSDM 0 272 368 582
<< end >>
