magic
tech sky130A
magscale 1 2
timestamp 1739872317
<< nwell >>
rect -38 262 682 582
<< pwell >>
rect 0 28 644 204
rect 0 22 460 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 338 298 368 496
rect 424 298 454 496
rect 510 298 540 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 252 48 282 178
rect 338 48 368 178
rect 424 48 454 178
rect 510 48 540 178
<< ndiff >>
rect 27 150 80 178
rect 27 60 35 150
rect 69 60 80 150
rect 27 48 80 60
rect 110 48 166 178
rect 196 148 252 178
rect 196 72 207 148
rect 241 72 252 148
rect 196 48 252 72
rect 282 48 338 178
rect 368 90 424 178
rect 368 56 379 90
rect 413 56 424 90
rect 368 48 424 56
rect 454 150 510 178
rect 454 72 465 150
rect 499 72 510 150
rect 454 48 510 72
rect 540 148 617 178
rect 540 56 553 148
rect 587 56 617 148
rect 540 48 617 56
<< pdiff >>
rect 27 476 80 496
rect 27 368 35 476
rect 69 368 80 476
rect 27 298 80 368
rect 110 484 166 496
rect 110 436 121 484
rect 155 436 166 484
rect 110 298 166 436
rect 196 476 252 496
rect 196 352 207 476
rect 241 352 252 476
rect 196 298 252 352
rect 282 488 338 496
rect 282 436 293 488
rect 327 436 338 488
rect 282 298 338 436
rect 368 476 424 496
rect 368 368 379 476
rect 413 368 424 476
rect 368 298 424 368
rect 454 408 510 496
rect 454 306 465 408
rect 499 306 510 408
rect 454 298 510 306
rect 540 476 617 496
rect 540 368 551 476
rect 585 368 617 476
rect 540 298 617 368
<< ndiffc >>
rect 35 60 69 150
rect 207 72 241 148
rect 379 56 413 90
rect 465 72 499 150
rect 553 56 587 148
<< pdiffc >>
rect 35 368 69 476
rect 121 436 155 484
rect 207 352 241 476
rect 293 436 327 488
rect 379 368 413 476
rect 465 306 499 408
rect 551 368 585 476
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 424 496 454 522
rect 510 496 540 522
rect 80 266 110 298
rect 60 250 114 266
rect 60 216 70 250
rect 104 216 114 250
rect 60 200 114 216
rect 166 260 196 298
rect 252 260 282 298
rect 338 266 368 298
rect 166 250 282 260
rect 166 216 182 250
rect 216 216 282 250
rect 166 204 282 216
rect 80 178 110 200
rect 166 178 196 204
rect 252 178 282 204
rect 324 250 378 266
rect 324 216 334 250
rect 368 216 378 250
rect 324 200 378 216
rect 424 260 454 298
rect 510 266 540 298
rect 510 260 578 266
rect 424 250 578 260
rect 424 216 534 250
rect 568 216 578 250
rect 424 204 578 216
rect 338 178 368 200
rect 424 178 454 204
rect 510 200 578 204
rect 510 178 540 200
rect 80 22 110 48
rect 166 22 196 48
rect 252 22 282 48
rect 338 22 368 48
rect 424 22 454 48
rect 510 22 540 48
<< polycont >>
rect 70 216 104 250
rect 182 216 216 250
rect 334 216 368 250
rect 534 216 568 250
<< locali >>
rect 0 561 644 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 526 644 527
rect 35 476 69 492
rect 121 484 155 526
rect 121 420 155 436
rect 207 476 241 492
rect 69 368 207 386
rect 35 352 207 368
rect 293 488 327 526
rect 293 420 327 436
rect 379 476 585 492
rect 241 368 379 386
rect 413 458 551 476
rect 241 352 413 368
rect 465 408 499 424
rect 76 284 358 318
rect 76 266 110 284
rect 60 250 110 266
rect 324 266 358 284
rect 452 306 465 316
rect 551 352 585 368
rect 324 250 378 266
rect 60 216 70 250
rect 104 216 110 250
rect 60 200 110 216
rect 166 216 182 250
rect 216 216 282 250
rect 166 200 282 216
rect 324 216 334 250
rect 368 216 378 250
rect 324 200 378 216
rect 452 166 499 306
rect 534 250 584 318
rect 568 216 584 250
rect 534 198 584 216
rect 35 150 69 166
rect 35 21 69 60
rect 207 150 499 166
rect 207 148 465 150
rect 241 132 465 148
rect 207 56 241 72
rect 362 90 430 98
rect 362 56 379 90
rect 413 56 430 90
rect 465 56 499 72
rect 553 148 587 164
rect 379 21 413 56
rect 553 21 587 56
rect 0 17 644 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel comment s 0 0 0 0 4 aoi21_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 68 221 102 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 85 238 85 238 0 FreeSans 200 0 0 0 A
flabel locali s 187 204 221 238 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 204 221 204 221 0 FreeSans 200 0 0 0 B
flabel locali s 544 204 578 238 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 561 221 561 221 0 FreeSans 200 0 0 0 C
flabel locali s 459 204 493 238 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 476 221 476 221 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__aoi21_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 644 220
string MASKHINTS_NSDM 0 -38 644 209
string MASKHINTS_PSDM 0 273 644 582
<< end >>
