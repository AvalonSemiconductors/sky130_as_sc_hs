magic
tech sky130A
magscale 1 2
timestamp 1733678203
<< nwell >>
rect -38 262 314 582
<< pwell >>
rect 2 44 274 204
rect 26 -15 76 44
rect 26 -20 66 -15
<< locali >>
rect 0 526 8 562
rect 268 526 276 562
rect 0 -15 8 21
rect 268 -15 276 21
<< viali >>
rect 8 526 268 562
rect 8 -15 268 21
<< metal1 >>
rect 0 562 276 592
rect 0 526 8 562
rect 268 526 276 562
rect 0 496 276 526
rect 0 21 276 48
rect 0 -15 8 21
rect 268 -15 276 21
rect 0 -48 276 -15
<< labels >>
rlabel comment s 0 0 0 0 4 aaaaaa
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 0 496 276 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 0 -48 276 48 1 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
