magic
tech sky130A
magscale 1 2
timestamp 1749431900
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 0 22 460 204
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 264 298 294 496
rect 350 298 380 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 264 48 294 178
rect 350 48 380 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 140 166 178
rect 110 106 121 140
rect 155 106 166 140
rect 110 48 166 106
rect 196 95 264 178
rect 196 61 207 95
rect 241 61 264 95
rect 196 48 264 61
rect 294 134 350 178
rect 294 100 305 134
rect 339 100 350 134
rect 294 48 350 100
rect 380 95 433 178
rect 380 61 391 95
rect 425 61 433 95
rect 380 48 433 61
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 298 80 336
rect 110 298 166 496
rect 196 488 264 496
rect 196 406 207 488
rect 241 406 264 488
rect 196 298 264 406
rect 294 440 350 496
rect 294 406 305 440
rect 339 406 350 440
rect 294 298 350 406
rect 380 484 433 496
rect 380 450 391 484
rect 425 450 433 484
rect 380 298 433 450
<< ndiffc >>
rect 35 72 69 150
rect 121 106 155 140
rect 207 61 241 95
rect 305 100 339 134
rect 391 61 425 95
<< pdiffc >>
rect 35 336 69 476
rect 207 406 241 488
rect 305 406 339 440
rect 391 450 425 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 264 496 294 522
rect 350 496 380 522
rect 80 266 110 298
rect 166 266 196 298
rect 264 266 294 298
rect 350 266 380 298
rect 36 250 110 266
rect 36 216 46 250
rect 80 216 110 250
rect 36 200 110 216
rect 156 250 212 266
rect 156 216 168 250
rect 202 216 212 250
rect 156 200 212 216
rect 264 250 380 266
rect 264 216 276 250
rect 310 216 380 250
rect 264 200 380 216
rect 80 178 110 200
rect 166 178 196 200
rect 264 178 294 200
rect 350 178 380 200
rect 80 22 110 48
rect 166 22 196 48
rect 264 22 294 48
rect 350 22 380 48
<< polycont >>
rect 46 216 80 250
rect 168 216 202 250
rect 276 216 310 250
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 35 476 69 492
rect 207 488 241 526
rect 375 484 442 526
rect 207 390 241 406
rect 305 440 339 456
rect 375 450 391 484
rect 425 450 442 484
rect 339 406 394 416
rect 305 390 394 406
rect 312 382 394 390
rect 69 336 290 356
rect 35 322 290 336
rect 35 320 106 322
rect 34 250 80 286
rect 34 216 46 250
rect 34 200 80 216
rect 152 250 202 288
rect 256 280 290 322
rect 152 216 168 250
rect 152 198 202 216
rect 237 266 290 280
rect 237 250 310 266
rect 237 216 276 250
rect 237 200 310 216
rect 35 150 69 166
rect 237 164 271 200
rect 344 172 394 382
rect 340 166 394 172
rect 112 140 271 164
rect 112 106 121 140
rect 155 130 271 140
rect 305 154 394 166
rect 305 134 374 154
rect 112 90 155 106
rect 339 132 374 134
rect 35 21 69 72
rect 191 61 207 95
rect 241 61 257 95
rect 305 84 339 100
rect 375 95 442 98
rect 375 61 391 95
rect 425 61 442 95
rect 207 21 241 61
rect 375 60 442 61
rect 391 21 425 60
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
flabel locali 153 238 187 272 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 170 255 170 255 0 FreeSans 200 0 0 0 B
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__or2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 220
string MASKHINTS_NSDM 0 -38 460 209
string MASKHINTS_PSDM 0 273 460 582
<< end >>
