magic
tech sky130A
magscale 1 2
timestamp 1740360520
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 0 -4 460 204
rect 26 -20 90 -4
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 338 298 368 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 252 48 282 178
rect 338 48 368 178
<< ndiff >>
rect 27 156 80 178
rect 27 64 35 156
rect 69 64 80 156
rect 27 48 80 64
rect 110 154 166 178
rect 110 120 121 154
rect 155 120 166 154
rect 110 48 166 120
rect 196 92 252 178
rect 196 58 207 92
rect 241 58 252 92
rect 196 48 252 58
rect 282 150 338 178
rect 282 116 293 150
rect 327 116 338 150
rect 282 48 338 116
rect 368 92 433 178
rect 368 58 380 92
rect 414 58 433 92
rect 368 48 433 58
<< pdiff >>
rect 27 476 80 496
rect 27 344 35 476
rect 69 344 80 476
rect 27 298 80 344
rect 110 486 166 496
rect 110 410 121 486
rect 155 410 166 486
rect 110 298 166 410
rect 196 476 252 496
rect 196 340 207 476
rect 241 340 252 476
rect 196 298 252 340
rect 282 356 338 496
rect 282 322 293 356
rect 327 322 338 356
rect 282 298 338 322
rect 368 476 433 496
rect 368 442 386 476
rect 420 442 433 476
rect 368 298 433 442
<< ndiffc >>
rect 35 64 69 156
rect 121 120 155 154
rect 207 58 241 92
rect 293 116 327 150
rect 380 58 414 92
<< pdiffc >>
rect 35 344 69 476
rect 121 410 155 486
rect 207 340 241 476
rect 293 322 327 356
rect 386 442 420 476
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 80 268 110 298
rect 166 268 196 298
rect 252 268 282 298
rect 338 268 368 298
rect 62 250 196 268
rect 62 216 94 250
rect 180 216 196 250
rect 62 200 196 216
rect 238 250 370 268
rect 238 216 254 250
rect 306 216 370 250
rect 238 200 370 216
rect 80 178 110 200
rect 166 178 196 200
rect 252 178 282 200
rect 338 178 368 200
rect 80 22 110 48
rect 166 22 196 48
rect 252 22 282 48
rect 338 22 368 48
<< polycont >>
rect 94 216 180 250
rect 254 216 306 250
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 34 476 70 492
rect 34 344 35 476
rect 69 348 70 476
rect 110 486 166 526
rect 110 410 121 486
rect 155 410 166 486
rect 110 394 166 410
rect 206 476 420 492
rect 206 348 207 476
rect 69 344 207 348
rect 34 340 207 344
rect 241 458 386 476
rect 241 340 242 458
rect 386 426 420 442
rect 34 314 242 340
rect 292 356 328 372
rect 292 322 293 356
rect 327 350 328 356
rect 327 322 432 350
rect 292 304 432 322
rect 78 250 196 268
rect 78 216 94 250
rect 180 216 196 250
rect 78 212 196 216
rect 238 250 322 268
rect 238 216 254 250
rect 306 216 322 250
rect 238 212 322 216
rect 374 178 432 304
rect 35 156 69 172
rect 120 154 432 178
rect 120 120 121 154
rect 155 150 432 154
rect 155 142 293 150
rect 155 120 156 142
rect 120 104 156 120
rect 292 116 293 142
rect 327 142 432 150
rect 327 116 328 142
rect 35 21 69 64
rect 207 92 241 108
rect 292 100 328 116
rect 207 21 241 58
rect 380 92 414 108
rect 380 21 414 58
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nor2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 A
flabel locali 255 221 289 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 272 238 272 238 0 FreeSans 200 0 0 0 B
flabel locali 391 187 425 221 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 408 204 408 204 0 FreeSans 200 0 0 0 Y
flabel locali 391 289 425 323 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 408 306 408 306 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__nor2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 214
string MASKHINTS_NSDM 0 -38 460 203
string MASKHINTS_PSDM 0 273 460 582
<< end >>
