magic
tech sky130A
magscale 1 2
timestamp 1739729400
<< nwell >>
rect -38 262 866 582
<< pwell >>
rect 22 48 820 204
rect 26 44 320 48
rect 26 24 90 44
rect 26 22 110 24
rect 26 -20 90 22
<< pmos >>
rect 80 375 110 496
rect 176 375 206 496
rect 266 375 296 496
rect 416 393 446 496
rect 512 393 542 496
rect 632 339 662 496
rect 718 339 748 496
<< nmoslvt >>
rect 80 48 110 138
rect 176 48 206 138
rect 266 48 296 138
rect 382 48 412 138
rect 512 48 542 168
rect 632 48 662 178
rect 718 48 748 178
<< ndiff >>
rect 586 168 632 178
rect 452 138 512 168
rect 27 114 80 138
rect 27 74 35 114
rect 69 74 80 114
rect 27 48 80 74
rect 110 102 176 138
rect 110 64 121 102
rect 155 64 176 102
rect 110 48 176 64
rect 206 48 266 138
rect 296 108 382 138
rect 296 74 308 108
rect 370 74 382 108
rect 296 48 382 74
rect 412 48 512 138
rect 542 92 632 168
rect 542 58 587 92
rect 621 58 632 92
rect 542 48 632 58
rect 662 170 718 178
rect 662 72 673 170
rect 707 72 718 170
rect 662 48 718 72
rect 748 166 801 178
rect 748 62 759 166
rect 793 62 801 166
rect 748 48 801 62
<< pdiff >>
rect 27 472 80 496
rect 27 410 35 472
rect 69 410 80 472
rect 27 375 80 410
rect 110 488 176 496
rect 110 452 121 488
rect 155 452 176 488
rect 110 375 176 452
rect 206 375 266 496
rect 296 474 416 496
rect 296 418 330 474
rect 382 418 416 474
rect 296 393 416 418
rect 446 393 512 496
rect 542 488 632 496
rect 542 404 574 488
rect 621 404 632 488
rect 542 393 632 404
rect 296 375 349 393
rect 582 339 632 393
rect 662 466 718 496
rect 662 350 673 466
rect 707 350 718 466
rect 662 339 718 350
rect 748 484 801 496
rect 748 388 759 484
rect 793 388 801 484
rect 748 339 801 388
<< ndiffc >>
rect 35 74 69 114
rect 121 64 155 102
rect 308 74 370 108
rect 587 58 621 92
rect 673 72 707 170
rect 759 62 793 166
<< pdiffc >>
rect 35 410 69 472
rect 121 452 155 488
rect 330 418 382 474
rect 574 404 621 488
rect 673 350 707 466
rect 759 388 793 484
<< poly >>
rect 80 496 110 522
rect 176 496 206 522
rect 266 496 296 522
rect 416 496 446 522
rect 512 496 542 522
rect 632 496 662 522
rect 718 496 748 522
rect 80 228 110 375
rect 176 334 206 375
rect 266 344 296 375
rect 416 362 446 393
rect 416 346 470 362
rect 152 318 206 334
rect 152 284 162 318
rect 196 284 206 318
rect 152 266 206 284
rect 248 328 306 344
rect 248 294 258 328
rect 292 298 306 328
rect 416 312 426 346
rect 460 312 470 346
rect 292 294 374 298
rect 416 296 470 312
rect 248 268 374 294
rect 80 212 134 228
rect 80 178 90 212
rect 124 178 134 212
rect 80 162 134 178
rect 80 138 110 162
rect 176 138 206 266
rect 248 210 302 226
rect 248 176 258 210
rect 292 176 302 210
rect 248 160 302 176
rect 344 194 374 268
rect 512 254 542 393
rect 632 308 662 339
rect 464 244 542 254
rect 464 210 484 244
rect 518 210 542 244
rect 588 302 662 308
rect 718 302 748 339
rect 588 292 748 302
rect 588 258 598 292
rect 632 258 748 292
rect 588 242 748 258
rect 464 198 542 210
rect 344 164 412 194
rect 512 168 542 198
rect 632 208 748 242
rect 632 178 662 208
rect 718 178 748 208
rect 266 138 296 160
rect 382 138 412 164
rect 80 22 110 48
rect 176 22 206 48
rect 266 22 296 48
rect 382 22 412 48
rect 512 22 542 48
rect 632 22 662 48
rect 718 22 748 48
<< polycont >>
rect 162 284 196 318
rect 258 294 292 328
rect 426 312 460 346
rect 90 178 124 212
rect 258 176 292 210
rect 484 210 518 244
rect 598 258 632 292
<< locali >>
rect 0 561 828 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 526 828 527
rect 121 488 155 526
rect 22 472 69 488
rect 22 410 35 472
rect 574 488 626 526
rect 121 436 155 452
rect 314 474 398 476
rect 22 402 69 410
rect 314 418 330 474
rect 382 430 398 474
rect 382 418 540 430
rect 22 368 274 402
rect 314 396 540 418
rect 22 132 56 368
rect 240 344 274 368
rect 416 350 470 362
rect 344 346 470 350
rect 90 318 206 334
rect 90 284 162 318
rect 196 284 206 318
rect 90 268 206 284
rect 240 328 292 344
rect 240 294 258 328
rect 240 278 292 294
rect 344 312 426 346
rect 460 312 470 346
rect 506 346 540 396
rect 621 404 626 488
rect 574 388 626 404
rect 673 466 707 486
rect 759 484 793 526
rect 759 372 793 388
rect 506 312 630 346
rect 344 296 470 312
rect 572 308 630 312
rect 673 338 707 350
rect 90 226 136 228
rect 90 224 298 226
rect 344 224 384 296
rect 572 292 639 308
rect 90 212 384 224
rect 124 210 384 212
rect 124 178 258 210
rect 90 176 258 178
rect 292 180 384 210
rect 440 244 538 262
rect 440 210 484 244
rect 518 210 538 244
rect 572 258 598 292
rect 632 258 639 292
rect 572 242 639 258
rect 292 176 298 180
rect 90 162 298 176
rect 248 160 298 162
rect 440 158 480 210
rect 572 176 606 242
rect 516 142 606 176
rect 673 224 748 338
rect 673 170 707 224
rect 22 114 69 132
rect 516 124 550 142
rect 22 100 35 114
rect 35 58 69 74
rect 121 102 155 118
rect 121 21 155 64
rect 296 108 550 124
rect 296 74 308 108
rect 370 90 550 108
rect 584 92 628 108
rect 370 74 384 90
rect 296 58 384 74
rect 584 58 587 92
rect 621 58 628 92
rect 584 21 628 58
rect 673 56 707 72
rect 759 166 793 188
rect 759 21 793 62
rect 0 17 828 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 170 170 204 204 0 FreeSans 200 0 0 0 S
port 8 nsew signal input
flabel locali 187 187 187 187 0 FreeSans 200 0 0 0 S
flabel locali 153 289 187 323 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 170 306 170 306 0 FreeSans 200 0 0 0 B
flabel locali 442 221 476 255 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel locali 459 238 459 238 0 FreeSans 200 0 0 0 A
flabel locali 697 255 731 289 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali 714 272 714 272 0 FreeSans 200 0 0 0 Y
flabel locali 425 306 459 340 0 FreeSans 200 0 0 0 S
port 8 nsew signal input
flabel locali 442 323 442 323 0 FreeSans 200 0 0 0 S
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__mux2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 828 216
string MASKHINTS_NSDM 0 -34 828 204
string MASKHINTS_PSDM 0 289 828 578
<< end >>
