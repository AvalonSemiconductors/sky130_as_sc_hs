magic
tech sky130A
magscale 1 2
timestamp 1733768868
<< nwell >>
rect -38 262 406 582
<< pwell >>
rect 24 44 320 204
rect 24 -15 76 44
rect 24 -22 70 -15
<< nmos >>
rect 118 56 158 194
rect 218 56 258 194
<< pmos >>
rect 118 322 158 496
rect 218 322 258 496
<< ndiff >>
rect 54 174 118 194
rect 54 66 70 174
rect 104 66 118 174
rect 54 56 118 66
rect 158 186 218 194
rect 158 80 172 186
rect 206 80 218 186
rect 158 56 218 80
rect 258 172 312 194
rect 258 68 270 172
rect 304 68 312 172
rect 258 56 312 68
<< pdiff >>
rect 56 488 118 496
rect 56 344 70 488
rect 104 344 118 488
rect 56 322 118 344
rect 158 460 218 496
rect 158 330 172 460
rect 206 330 218 460
rect 158 322 218 330
rect 258 488 318 496
rect 258 344 270 488
rect 304 344 318 488
rect 258 322 318 344
<< ndiffc >>
rect 70 66 104 174
rect 172 80 206 186
rect 270 68 304 172
<< pdiffc >>
rect 70 344 104 488
rect 172 330 206 460
rect 270 344 304 488
<< poly >>
rect 118 496 158 522
rect 218 496 258 522
rect 118 288 158 322
rect 60 272 158 288
rect 218 272 258 322
rect 60 238 76 272
rect 110 238 258 272
rect 60 232 258 238
rect 60 224 158 232
rect 118 194 158 224
rect 218 194 258 232
rect 118 30 158 56
rect 218 30 258 56
<< polycont >>
rect 76 238 110 272
<< locali >>
rect 0 561 368 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 526 368 527
rect 64 488 114 526
rect 64 344 70 488
rect 104 344 114 488
rect 264 488 314 526
rect 64 322 114 344
rect 164 460 214 486
rect 164 330 172 460
rect 206 330 214 460
rect 60 272 126 288
rect 60 238 76 272
rect 110 238 126 272
rect 60 224 126 238
rect 62 174 112 190
rect 62 66 70 174
rect 104 66 112 174
rect 62 21 112 66
rect 164 186 214 330
rect 264 344 270 488
rect 304 344 314 488
rect 264 322 314 344
rect 164 80 172 186
rect 206 80 214 186
rect 164 62 214 80
rect 256 172 310 190
rect 256 68 270 172
rect 304 68 310 172
rect 256 56 310 68
rect 256 21 306 56
rect 0 17 368 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -48 368 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 0 496 368 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 68 238 102 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 85 255 102 272 0 FreeSans 200 0 0 0 A
flabel locali 170 238 204 272 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 187 255 187 255 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__inv_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
