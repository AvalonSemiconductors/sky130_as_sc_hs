magic
tech sky130A
magscale 1 2
timestamp 1739791795
<< nwell >>
rect -38 262 1050 582
<< pwell >>
rect 0 26 1012 204
rect 0 24 920 26
rect 0 22 736 24
rect 782 22 812 24
rect 887 22 917 24
rect 26 -20 90 22
<< pmos >>
rect 80 347 110 496
rect 166 347 196 496
rect 284 298 314 496
rect 434 298 464 496
rect 672 298 702 496
rect 782 298 812 496
rect 887 298 917 496
<< nmoslvt >>
rect 80 48 110 166
rect 176 48 206 166
rect 284 48 314 178
rect 544 48 574 178
rect 672 48 702 178
rect 782 48 812 178
rect 887 48 917 178
<< ndiff >>
rect 230 166 284 178
rect 27 154 80 166
rect 27 72 35 154
rect 69 72 80 154
rect 27 48 80 72
rect 110 102 176 166
rect 110 68 121 102
rect 155 68 176 102
rect 110 48 176 68
rect 206 48 284 166
rect 314 150 544 178
rect 314 72 329 150
rect 363 90 544 150
rect 363 72 398 90
rect 314 56 398 72
rect 432 56 544 90
rect 314 48 544 56
rect 574 170 672 178
rect 574 72 624 170
rect 658 72 672 170
rect 574 48 672 72
rect 702 150 782 178
rect 702 58 718 150
rect 752 58 782 150
rect 702 48 782 58
rect 812 150 887 178
rect 812 72 842 150
rect 876 72 887 150
rect 812 48 887 72
rect 917 134 984 178
rect 917 58 928 134
rect 962 58 984 134
rect 917 48 984 58
<< pdiff >>
rect 27 472 80 496
rect 27 438 35 472
rect 69 438 80 472
rect 27 347 80 438
rect 110 474 166 496
rect 110 440 121 474
rect 155 440 166 474
rect 110 347 166 440
rect 196 347 284 496
rect 230 298 284 347
rect 314 466 434 496
rect 314 432 329 466
rect 363 432 434 466
rect 314 298 434 432
rect 464 346 672 496
rect 464 312 488 346
rect 522 312 564 346
rect 598 312 672 346
rect 464 298 672 312
rect 702 488 782 496
rect 702 454 716 488
rect 750 454 782 488
rect 702 298 782 454
rect 812 470 887 496
rect 812 322 842 470
rect 876 322 887 470
rect 812 298 887 322
rect 917 488 984 496
rect 917 338 938 488
rect 972 338 984 488
rect 917 298 984 338
<< ndiffc >>
rect 35 72 69 154
rect 121 68 155 102
rect 329 72 363 150
rect 398 56 432 90
rect 624 72 658 170
rect 718 58 752 150
rect 842 72 876 150
rect 928 58 962 134
<< pdiffc >>
rect 35 438 69 472
rect 121 440 155 474
rect 329 432 363 466
rect 488 312 522 346
rect 564 312 598 346
rect 716 454 750 488
rect 842 322 876 470
rect 938 338 972 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 284 496 314 522
rect 434 496 464 522
rect 672 496 702 522
rect 782 496 812 522
rect 887 496 917 522
rect 80 332 110 347
rect 166 332 196 347
rect 80 302 196 332
rect 80 296 133 302
rect 79 280 133 296
rect 79 246 89 280
rect 123 246 133 280
rect 284 266 314 298
rect 79 230 133 246
rect 176 250 242 260
rect 80 166 110 230
rect 176 216 192 250
rect 226 216 242 250
rect 176 206 242 216
rect 284 250 392 266
rect 284 216 346 250
rect 380 216 392 250
rect 176 166 206 206
rect 284 200 392 216
rect 434 260 464 298
rect 672 266 702 298
rect 782 266 812 298
rect 887 266 917 298
rect 434 250 502 260
rect 434 216 450 250
rect 484 216 502 250
rect 434 206 502 216
rect 544 250 598 266
rect 544 216 554 250
rect 588 216 598 250
rect 544 200 598 216
rect 672 250 740 266
rect 672 216 692 250
rect 726 216 740 250
rect 672 200 740 216
rect 782 250 917 266
rect 782 216 792 250
rect 826 216 917 250
rect 782 200 917 216
rect 284 178 314 200
rect 544 178 574 200
rect 672 178 702 200
rect 782 178 812 200
rect 887 178 917 200
rect 80 22 110 48
rect 176 22 206 48
rect 284 22 314 48
rect 544 22 574 48
rect 672 22 702 48
rect 782 22 812 48
rect 887 22 917 48
<< polycont >>
rect 89 246 123 280
rect 192 216 226 250
rect 346 216 380 250
rect 450 216 484 250
rect 554 216 588 250
rect 692 216 726 250
rect 792 216 826 250
<< locali >>
rect 0 561 1012 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 526 1012 527
rect 20 472 69 488
rect 20 418 35 472
rect 20 404 69 418
rect 121 474 155 526
rect 716 488 750 526
rect 329 466 363 488
rect 121 412 155 440
rect 278 432 329 446
rect 938 488 972 526
rect 363 432 682 446
rect 716 438 750 454
rect 842 470 876 486
rect 278 412 682 432
rect 20 186 55 404
rect 89 336 210 370
rect 89 280 140 336
rect 123 246 140 280
rect 89 220 140 246
rect 176 250 242 252
rect 176 216 192 250
rect 226 216 242 250
rect 176 208 242 216
rect 176 186 210 208
rect 20 154 210 186
rect 20 150 35 154
rect 69 152 210 154
rect 278 166 312 412
rect 648 402 682 412
rect 648 368 808 402
rect 472 334 488 346
rect 358 312 488 334
rect 522 312 564 346
rect 598 334 616 346
rect 598 312 658 334
rect 358 300 658 312
rect 358 266 392 300
rect 346 250 392 266
rect 380 216 392 250
rect 346 200 392 216
rect 434 250 502 260
rect 484 216 502 250
rect 434 214 502 216
rect 544 250 590 266
rect 544 216 554 250
rect 588 216 590 250
rect 544 200 590 216
rect 544 180 578 200
rect 426 166 578 180
rect 278 150 363 166
rect 278 128 329 150
rect 35 56 69 72
rect 121 102 155 118
rect 121 21 155 68
rect 460 146 578 166
rect 624 170 658 300
rect 774 266 808 368
rect 876 322 894 356
rect 938 322 972 338
rect 842 306 894 322
rect 860 300 894 306
rect 692 250 740 266
rect 726 216 740 250
rect 692 200 740 216
rect 774 250 826 266
rect 774 216 792 250
rect 774 200 826 216
rect 363 72 398 90
rect 329 56 398 72
rect 432 56 448 90
rect 860 180 912 300
rect 860 166 894 180
rect 624 56 658 72
rect 718 150 752 166
rect 718 21 752 58
rect 842 150 894 166
rect 876 130 894 150
rect 928 134 962 150
rect 842 56 876 72
rect 928 21 962 58
rect 0 17 1012 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 35 438 69 452
rect 35 418 69 438
rect 210 336 244 370
rect 434 216 450 250
rect 450 216 468 250
rect 426 132 460 166
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 22 454 80 458
rect 22 452 466 454
rect 22 418 35 452
rect 69 418 466 452
rect 22 416 466 418
rect 22 412 80 416
rect 198 370 282 382
rect 198 336 210 370
rect 244 336 282 370
rect 198 328 282 336
rect 248 182 282 328
rect 434 256 466 416
rect 422 250 480 256
rect 422 216 434 250
rect 468 216 480 250
rect 422 210 480 216
rect 248 166 472 182
rect 248 146 426 166
rect 414 132 426 146
rect 460 132 472 166
rect 414 126 472 132
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 102 238 136 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 697 221 731 255 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel locali 714 238 714 238 0 FreeSans 200 0 0 0 B
flabel polycont 119 255 119 255 0 FreeSans 200 0 0 0 A
flabel locali 867 221 901 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 881 238 881 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__xnor2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1012 214
string MASKHINTS_NSDM 0 -38 1012 204
string MASKHINTS_PSDM 0 272 1012 582
<< end >>
