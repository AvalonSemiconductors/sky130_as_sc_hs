magic
tech sky130A
magscale 1 2
timestamp 1734490064
<< nwell >>
rect -38 262 406 582
<< pwell >>
rect 6 42 362 204
rect 22 -20 90 42
<< pmos >>
rect 80 335 110 496
rect 168 335 198 496
rect 256 335 286 496
<< nmoslvt >>
rect 80 50 110 188
rect 168 50 198 188
rect 256 50 286 188
<< ndiff >>
rect 27 140 80 188
rect 27 76 35 140
rect 69 76 80 140
rect 27 50 80 76
rect 110 120 168 188
rect 110 58 121 120
rect 155 58 168 120
rect 110 50 168 58
rect 198 144 256 188
rect 198 74 210 144
rect 244 74 256 144
rect 198 50 256 74
rect 286 172 340 188
rect 286 64 298 172
rect 332 64 340 172
rect 286 50 340 64
<< pdiff >>
rect 27 466 80 496
rect 27 382 35 466
rect 69 382 80 466
rect 27 335 80 382
rect 110 488 168 496
rect 110 426 121 488
rect 155 426 168 488
rect 110 335 168 426
rect 198 468 256 496
rect 198 398 210 468
rect 244 398 256 468
rect 198 335 256 398
rect 286 482 340 496
rect 286 354 298 482
rect 332 354 340 482
rect 286 335 340 354
<< ndiffc >>
rect 35 76 69 140
rect 121 58 155 120
rect 210 74 244 144
rect 298 64 332 172
<< pdiffc >>
rect 35 382 69 466
rect 121 426 155 488
rect 210 398 244 468
rect 298 354 332 482
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 80 308 110 335
rect 28 288 110 308
rect 168 304 198 335
rect 28 254 44 288
rect 78 254 110 288
rect 28 238 110 254
rect 80 188 110 238
rect 152 288 206 304
rect 152 254 162 288
rect 196 282 206 288
rect 256 282 286 335
rect 196 254 286 282
rect 152 252 286 254
rect 152 242 206 252
rect 152 236 198 242
rect 168 188 198 236
rect 256 188 286 252
rect 80 24 110 50
rect 168 24 198 50
rect 256 24 286 50
<< polycont >>
rect 44 254 78 288
rect 162 254 196 288
<< locali >>
rect 0 561 368 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 526 368 527
rect 121 488 155 526
rect 35 466 69 484
rect 121 410 155 426
rect 210 468 264 484
rect 244 398 264 468
rect 210 382 264 398
rect 35 376 69 382
rect 35 342 176 376
rect 142 312 176 342
rect 31 288 90 308
rect 31 254 44 288
rect 78 254 90 288
rect 31 238 90 254
rect 142 288 196 312
rect 142 254 162 288
rect 142 236 196 254
rect 230 298 264 382
rect 298 482 332 526
rect 298 338 332 354
rect 230 246 278 298
rect 142 204 176 236
rect 35 170 176 204
rect 35 140 69 170
rect 230 160 264 246
rect 210 144 264 160
rect 35 58 69 76
rect 121 120 155 136
rect 244 74 264 144
rect 210 58 264 74
rect 298 172 332 188
rect 121 21 155 58
rect 298 21 332 64
rect 0 17 368 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 368 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali s 238 255 272 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 255 272 255 272 0 FreeSans 200 0 0 0 Y
flabel locali s 221 408 255 442 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 238 425 238 425 0 FreeSans 200 0 0 0 Y
flabel locali s 221 102 255 136 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 238 119 238 119 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
