magic
tech sky130A
magscale 1 2
timestamp 1739983972
<< nwell >>
rect -38 262 958 582
<< pwell >>
rect 0 28 920 204
rect 0 22 736 28
rect 26 -20 90 22
<< pmos >>
rect 82 298 112 496
rect 168 298 198 496
rect 254 298 284 496
rect 340 298 370 496
rect 530 298 560 496
rect 618 298 648 496
rect 706 298 736 496
rect 792 298 822 496
<< nmoslvt >>
rect 82 48 112 178
rect 168 48 198 178
rect 254 48 284 178
rect 340 48 370 178
rect 530 48 560 178
rect 618 48 648 178
rect 706 48 736 178
rect 792 48 822 178
<< ndiff >>
rect 27 152 82 178
rect 27 72 35 152
rect 69 72 82 152
rect 27 48 82 72
rect 112 168 168 178
rect 112 134 123 168
rect 157 134 168 168
rect 112 48 168 134
rect 198 90 254 178
rect 198 56 209 90
rect 243 56 254 90
rect 198 48 254 56
rect 284 168 340 178
rect 284 134 295 168
rect 329 134 340 168
rect 284 48 340 134
rect 370 90 530 178
rect 370 56 381 90
rect 498 56 530 90
rect 370 48 530 56
rect 560 94 618 178
rect 560 60 573 94
rect 607 60 618 94
rect 560 48 618 60
rect 648 150 706 178
rect 648 72 659 150
rect 693 72 706 150
rect 648 48 706 72
rect 736 94 792 178
rect 736 60 747 94
rect 781 60 792 94
rect 736 48 792 60
rect 822 164 893 178
rect 822 74 833 164
rect 867 74 893 164
rect 822 48 893 74
<< pdiff >>
rect 27 476 82 496
rect 27 356 37 476
rect 71 356 82 476
rect 27 298 82 356
rect 112 488 168 496
rect 112 454 123 488
rect 157 454 168 488
rect 112 298 168 454
rect 198 476 254 496
rect 198 356 209 476
rect 243 356 254 476
rect 198 298 254 356
rect 284 408 340 496
rect 284 320 295 408
rect 329 320 340 408
rect 284 298 340 320
rect 370 476 423 496
rect 370 404 381 476
rect 415 404 423 476
rect 370 298 423 404
rect 477 476 530 496
rect 477 404 485 476
rect 519 404 530 476
rect 477 298 530 404
rect 560 408 618 496
rect 560 320 573 408
rect 607 320 618 408
rect 560 298 618 320
rect 648 476 706 496
rect 648 336 661 476
rect 695 336 706 476
rect 648 298 706 336
rect 736 488 792 496
rect 736 404 747 488
rect 781 404 792 488
rect 736 298 792 404
rect 822 476 893 496
rect 822 336 833 476
rect 867 336 893 476
rect 822 298 893 336
<< ndiffc >>
rect 35 72 69 152
rect 123 134 157 168
rect 209 56 243 90
rect 295 134 329 168
rect 381 56 498 90
rect 573 60 607 94
rect 659 72 693 150
rect 747 60 781 94
rect 833 74 867 164
<< pdiffc >>
rect 37 356 71 476
rect 123 454 157 488
rect 209 356 243 476
rect 295 320 329 408
rect 381 404 415 476
rect 485 404 519 476
rect 573 320 607 408
rect 661 336 695 476
rect 747 404 781 488
rect 833 336 867 476
<< poly >>
rect 82 496 112 522
rect 168 496 198 522
rect 254 496 284 522
rect 340 496 370 522
rect 530 496 560 522
rect 618 496 648 522
rect 706 496 736 522
rect 792 496 822 522
rect 82 272 112 298
rect 168 272 198 298
rect 62 250 198 272
rect 62 216 78 250
rect 182 216 198 250
rect 62 204 198 216
rect 82 178 112 204
rect 168 178 198 204
rect 254 272 284 298
rect 340 272 370 298
rect 254 250 370 272
rect 254 216 270 250
rect 304 216 370 250
rect 254 204 370 216
rect 254 178 284 204
rect 340 178 370 204
rect 530 272 560 298
rect 618 272 648 298
rect 530 250 648 272
rect 530 216 576 250
rect 610 216 648 250
rect 530 204 648 216
rect 530 178 560 204
rect 618 178 648 204
rect 706 272 736 298
rect 792 272 822 298
rect 706 250 822 272
rect 706 216 740 250
rect 774 216 822 250
rect 706 204 822 216
rect 706 178 736 204
rect 792 178 822 204
rect 82 22 112 48
rect 168 22 198 48
rect 254 22 284 48
rect 340 22 370 48
rect 530 22 560 48
rect 618 22 648 48
rect 706 22 736 48
rect 792 22 822 48
<< polycont >>
rect 78 216 182 250
rect 270 216 304 250
rect 576 216 610 250
rect 740 216 774 250
<< locali >>
rect 0 561 920 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 526 920 527
rect 36 476 72 492
rect 36 356 37 476
rect 71 374 72 476
rect 123 488 157 526
rect 123 428 157 454
rect 209 476 415 492
rect 71 356 209 374
rect 243 458 381 476
rect 36 340 243 356
rect 295 408 329 424
rect 278 320 295 354
rect 381 388 415 404
rect 485 476 695 492
rect 519 458 661 476
rect 485 388 519 404
rect 573 408 607 424
rect 329 320 573 354
rect 607 320 624 354
rect 747 488 781 526
rect 747 388 781 404
rect 833 476 867 492
rect 695 336 833 354
rect 661 320 867 336
rect 62 272 130 306
rect 62 250 198 272
rect 62 216 78 250
rect 182 216 198 250
rect 62 204 198 216
rect 232 250 324 272
rect 232 216 270 250
rect 304 216 324 250
rect 232 204 324 216
rect 358 168 432 320
rect 530 250 644 272
rect 530 216 576 250
rect 610 216 644 250
rect 530 204 644 216
rect 706 250 804 272
rect 706 216 740 250
rect 774 216 804 250
rect 706 204 804 216
rect 35 152 69 168
rect 104 134 123 168
rect 157 134 295 168
rect 329 134 432 168
rect 833 166 867 180
rect 482 164 867 166
rect 482 150 833 164
rect 482 132 659 150
rect 482 90 516 132
rect 69 72 209 90
rect 35 56 209 72
rect 243 56 381 90
rect 498 56 516 90
rect 554 94 624 98
rect 554 60 573 94
rect 607 60 624 94
rect 693 132 833 150
rect 573 21 607 60
rect 659 56 693 72
rect 728 94 799 98
rect 728 60 747 94
rect 781 60 799 94
rect 747 21 781 60
rect 833 58 867 74
rect 0 17 920 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 oai22_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 68 221 102 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 85 238 85 238 0 FreeSans 200 0 0 0 A
flabel locali s 238 221 272 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 255 238 255 238 0 FreeSans 200 0 0 0 B
flabel locali s 561 221 595 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 578 238 578 238 0 FreeSans 200 0 0 0 C
flabel locali s 731 221 765 255 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel locali s 748 238 748 238 0 FreeSans 200 0 0 0 D
flabel locali s 391 221 425 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 408 238 408 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__oai22_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 920 220
string MASKHINTS_NSDM 0 -38 920 209
string MASKHINTS_PSDM 0 273 920 582
<< end >>
