magic
tech sky130A
magscale 1 2
timestamp 1740839465
<< nwell >>
rect -38 262 956 582
<< pwell >>
rect 0 32 920 204
rect 0 24 918 32
rect 0 22 736 24
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 186 298 216 496
rect 388 298 418 496
rect 474 298 504 496
rect 570 298 600 496
rect 664 298 694 496
rect 782 298 812 496
<< nmoslvt >>
rect 80 48 110 178
rect 186 48 216 178
rect 276 48 306 178
rect 380 48 410 178
rect 570 48 600 178
rect 682 48 712 178
rect 782 48 812 178
<< ndiff >>
rect 27 142 80 178
rect 27 108 35 142
rect 69 108 80 142
rect 27 48 80 108
rect 110 90 186 178
rect 110 56 121 90
rect 155 56 186 90
rect 110 48 186 56
rect 216 48 276 178
rect 306 96 380 178
rect 306 62 324 96
rect 358 62 380 96
rect 306 48 380 62
rect 410 48 570 178
rect 600 94 682 178
rect 600 60 628 94
rect 662 60 682 94
rect 600 48 682 60
rect 712 170 782 178
rect 712 136 737 170
rect 771 136 782 170
rect 712 48 782 136
rect 812 168 880 178
rect 812 56 823 168
rect 857 56 880 168
rect 812 48 880 56
<< pdiff >>
rect 27 476 80 496
rect 27 310 35 476
rect 69 310 80 476
rect 27 298 80 310
rect 110 488 186 496
rect 110 454 130 488
rect 164 454 186 488
rect 110 298 186 454
rect 216 298 388 496
rect 418 468 474 496
rect 418 434 429 468
rect 463 434 474 468
rect 418 298 474 434
rect 504 298 570 496
rect 600 484 664 496
rect 600 450 619 484
rect 653 450 664 484
rect 600 298 664 450
rect 694 476 782 496
rect 694 306 737 476
rect 771 306 782 476
rect 694 298 782 306
rect 812 488 880 496
rect 812 330 823 488
rect 857 330 880 488
rect 812 298 880 330
<< ndiffc >>
rect 35 108 69 142
rect 121 56 155 90
rect 324 62 358 96
rect 628 60 662 94
rect 737 136 771 170
rect 823 56 857 168
<< pdiffc >>
rect 35 310 69 476
rect 130 454 164 488
rect 429 434 463 468
rect 619 450 653 484
rect 737 306 771 476
rect 823 330 857 488
<< poly >>
rect 80 496 110 522
rect 186 496 216 522
rect 388 496 418 522
rect 474 496 504 522
rect 570 496 600 522
rect 664 496 694 522
rect 782 496 812 522
rect 80 266 110 298
rect 186 266 216 298
rect 388 266 418 298
rect 474 266 504 298
rect 570 266 600 298
rect 664 266 694 298
rect 80 250 136 266
rect 80 216 90 250
rect 124 216 136 250
rect 80 198 136 216
rect 178 250 232 266
rect 178 216 188 250
rect 222 216 232 250
rect 178 198 232 216
rect 274 250 328 266
rect 274 216 284 250
rect 318 216 328 250
rect 274 198 328 216
rect 370 250 424 266
rect 370 216 380 250
rect 414 216 424 250
rect 370 198 424 216
rect 466 250 520 266
rect 466 216 476 250
rect 510 216 520 250
rect 466 198 520 216
rect 562 250 616 266
rect 562 216 572 250
rect 606 216 616 250
rect 562 198 616 216
rect 658 250 712 266
rect 782 250 812 298
rect 658 216 668 250
rect 702 216 812 250
rect 658 198 712 216
rect 80 178 110 198
rect 186 178 216 198
rect 276 178 306 198
rect 380 178 410 198
rect 570 178 600 198
rect 682 178 712 198
rect 782 178 812 216
rect 80 22 110 48
rect 186 22 216 48
rect 276 22 306 48
rect 380 22 410 48
rect 570 22 600 48
rect 682 22 712 48
rect 782 22 812 48
<< polycont >>
rect 90 216 124 250
rect 188 216 222 250
rect 284 216 318 250
rect 380 216 414 250
rect 476 216 510 250
rect 572 216 606 250
rect 668 216 702 250
<< locali >>
rect 0 561 920 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 526 920 527
rect 35 476 69 492
rect 20 310 35 328
rect 130 488 164 526
rect 619 484 653 526
rect 130 434 164 454
rect 410 434 429 468
rect 463 434 536 468
rect 619 434 653 450
rect 737 476 771 492
rect 69 366 414 400
rect 20 294 69 310
rect 20 158 54 294
rect 90 250 144 266
rect 124 216 144 250
rect 90 198 144 216
rect 182 250 224 330
rect 182 216 188 250
rect 222 216 224 250
rect 182 198 224 216
rect 284 250 318 266
rect 110 164 144 198
rect 284 164 318 216
rect 380 250 414 366
rect 502 396 536 434
rect 502 362 702 396
rect 474 266 516 328
rect 576 266 616 328
rect 380 198 414 216
rect 466 250 518 266
rect 466 216 476 250
rect 510 216 518 250
rect 466 198 518 216
rect 562 250 616 266
rect 562 216 572 250
rect 606 216 616 250
rect 562 198 616 216
rect 668 250 702 362
rect 476 164 510 198
rect 20 142 70 158
rect 18 108 35 142
rect 69 108 70 142
rect 110 130 510 164
rect 668 162 702 216
rect 34 92 70 108
rect 544 128 702 162
rect 823 488 857 526
rect 823 314 857 330
rect 737 300 771 306
rect 737 212 792 300
rect 737 170 771 212
rect 544 96 578 128
rect 737 120 771 136
rect 823 168 857 184
rect 104 56 121 90
rect 155 56 172 90
rect 298 62 324 96
rect 358 62 578 96
rect 612 60 628 94
rect 662 60 680 94
rect 119 21 155 56
rect 626 21 662 60
rect 823 21 857 56
rect 0 17 920 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 mux2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 102 221 136 255 0 FreeSans 200 0 0 0 S
port 5 nsew signal input
flabel locali s 119 238 119 238 0 FreeSans 200 0 0 0 S
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 B
flabel locali s 476 221 510 255 0 FreeSans 200 0 0 0 S
port 5 nsew signal input
flabel locali s 493 238 493 238 0 FreeSans 200 0 0 0 S
flabel locali s 578 221 612 255 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel locali s 595 238 595 238 0 FreeSans 200 0 0 0 A
flabel locali s 748 221 782 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 765 238 765 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__mux2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 920 214
string MASKHINTS_NSDM 0 -38 920 204
string MASKHINTS_PSDM 0 272 920 582
<< end >>
