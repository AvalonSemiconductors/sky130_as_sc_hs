magic
tech sky130A
magscale 1 2
timestamp 1740561655
<< nwell >>
rect -38 262 590 582
<< pwell >>
rect 0 34 552 204
rect 0 22 460 34
rect 26 -20 90 22
<< pmos >>
rect 132 298 162 496
rect 226 298 256 496
rect 356 298 386 496
rect 442 298 472 496
<< nmoslvt >>
rect 132 48 162 178
rect 226 48 256 178
rect 356 48 386 178
rect 442 48 472 178
<< ndiff >>
rect 74 164 132 178
rect 74 130 87 164
rect 121 130 132 164
rect 74 48 132 130
rect 162 48 226 178
rect 256 94 356 178
rect 256 60 311 94
rect 345 60 356 94
rect 256 48 356 60
rect 386 170 442 178
rect 386 136 397 170
rect 431 136 442 170
rect 386 48 442 136
rect 472 166 525 178
rect 472 60 483 166
rect 517 60 525 166
rect 472 48 525 60
<< pdiff >>
rect 72 488 132 496
rect 72 316 85 488
rect 119 316 132 488
rect 72 298 132 316
rect 162 434 226 496
rect 162 328 176 434
rect 210 328 226 434
rect 162 298 226 328
rect 256 488 356 496
rect 256 420 286 488
rect 320 420 356 488
rect 256 298 356 420
rect 386 476 442 496
rect 386 306 397 476
rect 431 306 442 476
rect 386 298 442 306
rect 472 484 525 496
rect 472 338 483 484
rect 517 338 525 484
rect 472 298 525 338
<< ndiffc >>
rect 87 130 121 164
rect 311 60 345 94
rect 397 136 431 170
rect 483 60 517 166
<< pdiffc >>
rect 85 316 119 488
rect 176 328 210 434
rect 286 420 320 488
rect 397 306 431 476
rect 483 338 517 484
<< poly >>
rect 132 496 162 522
rect 226 496 256 522
rect 356 496 386 522
rect 442 496 472 522
rect 132 266 162 298
rect 226 266 256 298
rect 356 266 386 298
rect 116 250 170 266
rect 116 216 126 250
rect 160 216 170 250
rect 116 198 170 216
rect 222 250 276 266
rect 222 216 232 250
rect 266 216 276 250
rect 222 198 276 216
rect 318 264 386 266
rect 442 264 472 298
rect 318 250 472 264
rect 318 216 328 250
rect 362 216 472 250
rect 318 198 472 216
rect 132 178 162 198
rect 226 178 256 198
rect 356 178 386 198
rect 442 178 472 198
rect 132 22 162 48
rect 226 22 256 48
rect 356 22 386 48
rect 442 22 472 48
<< polycont >>
rect 126 216 160 250
rect 232 216 266 250
rect 328 216 362 250
<< locali >>
rect 0 561 552 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 526 552 527
rect 85 488 119 526
rect 286 488 320 526
rect 85 300 119 316
rect 176 434 210 450
rect 286 402 320 420
rect 397 476 431 492
rect 210 328 362 346
rect 176 312 362 328
rect 68 250 170 266
rect 68 216 126 250
rect 160 216 170 250
rect 68 198 170 216
rect 222 250 276 278
rect 222 216 232 250
rect 266 216 276 250
rect 222 198 276 216
rect 328 250 362 312
rect 328 164 362 216
rect 71 130 87 164
rect 121 130 362 164
rect 483 484 517 526
rect 483 322 517 338
rect 397 296 431 306
rect 397 214 460 296
rect 397 170 431 214
rect 397 120 431 136
rect 483 166 517 182
rect 294 94 362 96
rect 294 60 311 94
rect 345 60 362 94
rect 311 21 345 60
rect 483 21 517 60
rect 0 17 552 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 68 221 102 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 85 238 85 238 0 FreeSans 200 0 0 0 A
flabel locali s 238 221 272 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 255 238 255 238 0 FreeSans 200 0 0 0 B
flabel locali s 408 221 442 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 425 238 425 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__and2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 552 220
string MASKHINTS_NSDM 0 -38 552 209
string MASKHINTS_PSDM 0 273 552 582
<< end >>
