magic
tech sky130A
magscale 1 2
timestamp 1740921530
<< nwell >>
rect -38 262 682 582
<< pwell >>
rect 0 26 644 204
rect 0 22 460 26
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 268 298 298 496
rect 354 298 384 496
rect 440 298 470 496
rect 526 298 556 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 268 48 298 178
rect 354 48 384 178
rect 440 48 470 178
rect 526 48 556 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 140 166 178
rect 110 106 121 140
rect 155 106 166 140
rect 110 48 166 106
rect 196 150 268 178
rect 196 72 207 150
rect 241 72 268 150
rect 196 48 268 72
rect 298 140 354 178
rect 298 106 309 140
rect 343 106 354 140
rect 298 48 354 106
rect 384 95 440 178
rect 384 61 395 95
rect 429 61 440 95
rect 384 48 440 61
rect 470 170 526 178
rect 470 136 481 170
rect 515 136 526 170
rect 470 48 526 136
rect 556 166 609 178
rect 556 60 567 166
rect 601 60 609 166
rect 556 48 609 60
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 298 80 336
rect 110 298 166 496
rect 196 488 268 496
rect 196 406 207 488
rect 241 406 268 488
rect 196 298 268 406
rect 298 440 354 496
rect 298 406 309 440
rect 343 406 354 440
rect 298 298 354 406
rect 384 484 440 496
rect 384 450 395 484
rect 429 450 440 484
rect 384 298 440 450
rect 470 476 526 496
rect 470 306 481 476
rect 515 306 526 476
rect 470 298 526 306
rect 556 488 617 496
rect 556 306 567 488
rect 601 306 617 488
rect 556 298 617 306
<< ndiffc >>
rect 35 72 69 150
rect 121 106 155 140
rect 207 72 241 150
rect 309 106 343 140
rect 395 61 429 95
rect 481 136 515 170
rect 567 60 601 166
<< pdiffc >>
rect 35 336 69 476
rect 207 406 241 488
rect 309 406 343 440
rect 395 450 429 484
rect 481 306 515 476
rect 567 306 601 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 268 496 298 522
rect 354 496 384 522
rect 440 496 470 522
rect 526 496 556 522
rect 80 266 110 298
rect 36 250 110 266
rect 36 216 46 250
rect 80 216 110 250
rect 36 200 110 216
rect 80 178 110 200
rect 166 266 196 298
rect 268 266 298 298
rect 354 266 384 298
rect 166 250 226 266
rect 166 216 182 250
rect 216 216 226 250
rect 166 200 226 216
rect 268 250 384 266
rect 268 216 278 250
rect 312 244 384 250
rect 440 244 470 298
rect 312 238 470 244
rect 526 238 556 298
rect 312 216 556 238
rect 268 200 556 216
rect 166 178 196 200
rect 268 178 298 200
rect 354 178 384 200
rect 440 178 470 200
rect 526 178 556 200
rect 80 22 110 48
rect 166 22 196 48
rect 268 22 298 48
rect 354 22 384 48
rect 440 22 470 48
rect 526 22 556 48
<< polycont >>
rect 46 216 80 250
rect 182 216 216 250
rect 278 216 312 250
<< locali >>
rect 0 561 644 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 526 644 527
rect 35 476 69 492
rect 207 488 241 526
rect 378 484 446 526
rect 207 390 241 406
rect 303 440 343 456
rect 378 450 395 484
rect 429 450 446 484
rect 481 476 516 492
rect 303 406 309 440
rect 343 406 392 416
rect 303 390 392 406
rect 314 382 392 390
rect 69 348 292 356
rect 69 336 295 348
rect 35 322 295 336
rect 35 320 148 322
rect 34 250 80 286
rect 34 216 46 250
rect 34 200 80 216
rect 114 172 148 320
rect 182 250 226 288
rect 216 216 226 250
rect 182 200 226 216
rect 261 266 295 322
rect 261 250 312 266
rect 261 216 278 250
rect 261 200 312 216
rect 346 254 392 382
rect 515 306 516 476
rect 481 254 516 306
rect 567 488 601 526
rect 567 286 601 306
rect 346 220 516 254
rect 35 150 69 166
rect 114 140 155 172
rect 346 166 388 220
rect 114 106 121 140
rect 114 90 155 106
rect 207 150 241 166
rect 35 21 69 72
rect 303 154 388 166
rect 480 170 516 220
rect 303 140 380 154
rect 303 106 309 140
rect 343 132 380 140
rect 480 136 481 170
rect 515 136 516 170
rect 480 120 516 136
rect 567 166 601 182
rect 303 90 343 106
rect 378 95 446 98
rect 207 21 241 72
rect 378 61 395 95
rect 429 61 446 95
rect 378 60 446 61
rect 391 21 425 60
rect 567 21 601 60
rect 0 17 644 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 B
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__or2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 644 220
string MASKHINTS_NSDM 0 -38 644 209
string MASKHINTS_PSDM 0 273 644 582
<< end >>
