magic
tech sky130A
magscale 1 2
timestamp 1740359326
<< nwell >>
rect -38 262 682 582
<< pwell >>
rect 0 26 644 204
rect 0 22 460 26
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 262 298 292 496
rect 350 298 380 496
rect 436 298 466 496
rect 522 298 552 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 262 48 292 178
rect 350 48 380 178
rect 436 48 466 178
rect 522 48 552 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 140 166 178
rect 110 106 121 140
rect 155 106 166 140
rect 110 48 166 106
rect 196 150 262 178
rect 196 72 207 150
rect 241 72 262 150
rect 196 48 262 72
rect 292 140 350 178
rect 292 106 303 140
rect 337 106 350 140
rect 292 48 350 106
rect 380 95 436 178
rect 380 61 391 95
rect 425 61 436 95
rect 380 48 436 61
rect 466 170 522 178
rect 466 72 477 170
rect 511 72 522 170
rect 466 48 522 72
rect 552 166 607 178
rect 552 60 563 166
rect 597 60 607 166
rect 552 48 607 60
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 298 80 336
rect 110 298 166 496
rect 196 488 262 496
rect 196 406 207 488
rect 241 406 262 488
rect 196 298 262 406
rect 292 440 350 496
rect 292 406 303 440
rect 337 406 350 440
rect 292 298 350 406
rect 380 484 436 496
rect 380 450 391 484
rect 425 450 436 484
rect 380 298 436 450
rect 466 476 522 496
rect 466 306 477 476
rect 511 306 522 476
rect 466 298 522 306
rect 552 488 617 496
rect 552 306 563 488
rect 597 306 617 488
rect 552 298 617 306
<< ndiffc >>
rect 35 72 69 150
rect 121 106 155 140
rect 207 72 241 150
rect 303 106 337 140
rect 391 61 425 95
rect 477 72 511 170
rect 563 60 597 166
<< pdiffc >>
rect 35 336 69 476
rect 207 406 241 488
rect 303 406 337 440
rect 391 450 425 484
rect 477 306 511 476
rect 563 306 597 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 262 496 292 522
rect 350 496 380 522
rect 436 496 466 522
rect 522 496 552 522
rect 80 266 110 298
rect 30 250 110 266
rect 30 216 40 250
rect 74 216 110 250
rect 30 200 110 216
rect 80 178 110 200
rect 166 266 196 298
rect 262 266 292 298
rect 350 266 380 298
rect 166 250 220 266
rect 166 216 176 250
rect 210 216 220 250
rect 166 200 220 216
rect 262 250 380 266
rect 262 216 272 250
rect 306 244 380 250
rect 436 244 466 298
rect 306 238 466 244
rect 522 238 552 298
rect 306 216 552 238
rect 262 200 552 216
rect 166 178 196 200
rect 262 178 292 200
rect 350 178 380 200
rect 436 178 466 200
rect 522 178 552 200
rect 80 22 110 48
rect 166 22 196 48
rect 262 22 292 48
rect 350 22 380 48
rect 436 22 466 48
rect 522 22 552 48
<< polycont >>
rect 40 216 74 250
rect 176 216 210 250
rect 272 216 306 250
<< locali >>
rect 0 561 644 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 526 644 527
rect 35 476 69 492
rect 207 488 241 526
rect 374 484 442 526
rect 207 390 241 406
rect 303 440 337 456
rect 374 450 391 484
rect 425 450 442 484
rect 476 476 512 492
rect 337 406 392 416
rect 303 390 392 406
rect 312 382 392 390
rect 69 336 289 356
rect 35 322 289 336
rect 35 320 142 322
rect 30 250 74 286
rect 30 216 40 250
rect 30 200 74 216
rect 108 172 142 320
rect 176 250 221 288
rect 210 216 221 250
rect 176 200 221 216
rect 255 266 289 322
rect 255 250 306 266
rect 255 216 272 250
rect 255 200 306 216
rect 340 258 392 382
rect 476 306 477 476
rect 511 306 512 476
rect 340 254 400 258
rect 476 254 512 306
rect 563 488 597 526
rect 563 286 597 306
rect 340 220 512 254
rect 35 150 69 166
rect 108 140 155 172
rect 340 166 388 220
rect 108 106 121 140
rect 108 90 155 106
rect 207 150 241 166
rect 35 21 69 72
rect 303 154 388 166
rect 476 170 512 220
rect 303 140 374 154
rect 337 132 374 140
rect 303 90 337 106
rect 374 95 442 98
rect 207 21 241 72
rect 374 61 391 95
rect 425 61 442 95
rect 374 60 442 61
rect 476 72 477 170
rect 511 72 512 170
rect 391 21 425 60
rect 476 56 512 72
rect 563 166 597 182
rect 563 21 597 60
rect 0 17 644 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 187 221 221 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 204 238 204 238 0 FreeSans 200 0 0 0 B
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__or2_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 644 220
string MASKHINTS_NSDM 0 -38 644 209
string MASKHINTS_PSDM 0 273 644 582
<< end >>
