VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.605 2.050 0.775 2.630 ;
        RECT 1.490 1.690 1.660 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.680 ;
        RECT 1.490 0.105 1.660 0.940 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.210 1.810 1.020 ;
        RECT 0.110 -0.100 0.450 0.210 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.224250 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.190 0.450 1.540 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.433550 ;
    PORT
      LAYER li1 ;
        RECT 1.050 1.910 1.320 2.420 ;
        RECT 1.150 1.490 1.320 1.910 ;
        RECT 1.150 1.230 1.390 1.490 ;
        RECT 1.150 0.800 1.320 1.230 ;
        RECT 1.050 0.290 1.320 0.800 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.880 0.345 2.420 ;
        RECT 0.175 1.710 0.880 1.880 ;
        RECT 0.710 1.560 0.880 1.710 ;
        RECT 0.710 1.180 0.980 1.560 ;
        RECT 0.710 1.020 0.880 1.180 ;
        RECT 0.175 0.850 0.880 1.020 ;
        RECT 0.175 0.290 0.345 0.850 ;
  END
END sky130_as_sc_hs__buff_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__clkbuff_8
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__clkbuff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 5.260 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 5.070 2.810 ;
        RECT 0.130 1.540 0.400 2.630 ;
        RECT 1.000 1.850 1.270 2.630 ;
        RECT 1.880 1.850 2.150 2.630 ;
        RECT 2.780 1.850 3.050 2.630 ;
        RECT 3.660 1.850 3.930 2.630 ;
        RECT 4.540 1.850 4.810 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 5.070 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.105 0.390 0.670 ;
        RECT 1.010 0.105 1.260 0.550 ;
        RECT 1.890 0.105 2.140 0.550 ;
        RECT 2.790 0.105 3.040 0.560 ;
        RECT 3.670 0.105 3.920 0.560 ;
        RECT 4.550 0.105 4.800 0.560 ;
        RECT 0.000 -0.085 5.060 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 5.060 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.681500 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.680 1.710 2.460 ;
        RECT 2.390 1.680 2.610 2.460 ;
        RECT 3.220 1.680 3.490 2.460 ;
        RECT 4.100 1.680 4.370 2.460 ;
        RECT 1.490 1.510 4.910 1.680 ;
        RECT 4.050 0.900 4.910 1.510 ;
        RECT 1.490 0.730 4.910 0.900 ;
        RECT 1.490 0.280 1.700 0.730 ;
        RECT 2.390 0.280 2.600 0.730 ;
        RECT 3.230 0.280 3.480 0.730 ;
        RECT 4.110 0.280 4.360 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.427500 ;
    PORT
      LAYER li1 ;
        RECT 0.130 1.070 0.980 1.340 ;
        RECT 0.130 0.840 0.400 1.070 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.570 1.680 0.820 2.460 ;
        RECT 0.570 1.510 1.320 1.680 ;
        RECT 1.150 1.340 1.320 1.510 ;
        RECT 1.150 1.070 3.880 1.340 ;
        RECT 1.150 0.900 1.320 1.070 ;
        RECT 0.570 0.730 1.320 0.900 ;
        RECT 0.570 0.280 0.820 0.730 ;
  END
END sky130_as_sc_hs__clkbuff_8

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__buff_11
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__buff_11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.180 1.890 0.350 2.630 ;
        RECT 1.050 1.955 1.220 2.630 ;
        RECT 1.930 1.960 2.100 2.630 ;
        RECT 2.830 1.965 3.000 2.630 ;
        RECT 3.710 1.965 3.880 2.630 ;
        RECT 4.590 1.965 4.760 2.630 ;
        RECT 5.470 1.965 5.640 2.630 ;
        RECT 6.360 1.965 6.530 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.105 0.350 0.740 ;
        RECT 1.050 0.105 1.220 0.700 ;
        RECT 1.930 0.105 2.100 0.700 ;
        RECT 2.830 0.105 3.000 0.700 ;
        RECT 3.710 0.105 3.880 0.700 ;
        RECT 4.590 0.105 4.760 0.700 ;
        RECT 5.470 0.105 5.640 0.700 ;
        RECT 6.360 0.105 6.530 0.700 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 7.120 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.909000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 1.220 1.880 1.445 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.681550 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.795 2.560 2.460 ;
        RECT 3.270 1.795 3.440 2.460 ;
        RECT 4.150 1.795 4.320 2.460 ;
        RECT 5.030 1.795 5.200 2.460 ;
        RECT 5.920 1.795 6.090 2.460 ;
        RECT 6.800 1.795 6.970 2.460 ;
        RECT 2.390 1.625 7.220 1.795 ;
        RECT 6.890 1.040 7.220 1.625 ;
        RECT 2.390 0.870 7.220 1.040 ;
        RECT 2.390 0.280 2.560 0.870 ;
        RECT 3.270 0.280 3.440 0.870 ;
        RECT 4.150 0.280 4.320 0.870 ;
        RECT 5.030 0.280 5.200 0.870 ;
        RECT 5.910 0.280 6.080 0.870 ;
        RECT 6.800 0.280 6.970 0.870 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.610 1.785 0.780 2.460 ;
        RECT 1.490 1.785 1.660 2.460 ;
        RECT 0.610 1.615 2.220 1.785 ;
        RECT 2.050 1.455 2.220 1.615 ;
        RECT 2.050 1.230 6.720 1.455 ;
        RECT 2.050 1.050 2.220 1.230 ;
        RECT 0.610 0.870 2.220 1.050 ;
        RECT 0.610 0.280 0.780 0.870 ;
        RECT 1.490 0.280 1.660 0.870 ;
  END
END sky130_as_sc_hs__buff_11

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__clkbuff_11
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__clkbuff_11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.130 1.540 0.400 2.630 ;
        RECT 1.000 1.850 1.270 2.630 ;
        RECT 1.880 1.850 2.150 2.630 ;
        RECT 2.780 1.850 3.050 2.630 ;
        RECT 3.660 1.850 3.930 2.630 ;
        RECT 4.540 1.850 4.810 2.630 ;
        RECT 5.420 1.850 5.690 2.630 ;
        RECT 6.310 1.850 6.580 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.105 0.390 0.670 ;
        RECT 1.010 0.105 1.260 0.550 ;
        RECT 1.890 0.105 2.140 0.550 ;
        RECT 2.790 0.105 3.040 0.560 ;
        RECT 3.670 0.105 3.920 0.560 ;
        RECT 4.550 0.105 4.800 0.560 ;
        RECT 5.430 0.105 5.680 0.560 ;
        RECT 6.320 0.105 6.570 0.560 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.220 7.120 1.020 ;
        RECT 0.100 -0.075 0.410 0.220 ;
        RECT 0.100 -0.100 0.370 -0.075 ;
    END
  END VNB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.855000 ;
    PORT
      LAYER li1 ;
        RECT 0.260 1.070 1.870 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522250 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.680 2.610 2.460 ;
        RECT 3.220 1.680 3.490 2.460 ;
        RECT 4.100 1.680 4.370 2.460 ;
        RECT 4.980 1.680 5.250 2.460 ;
        RECT 5.870 1.680 6.140 2.460 ;
        RECT 6.750 1.870 7.020 2.460 ;
        RECT 6.750 1.680 7.200 1.870 ;
        RECT 2.390 1.510 7.200 1.680 ;
        RECT 6.690 0.900 7.200 1.510 ;
        RECT 2.390 0.730 7.200 0.900 ;
        RECT 2.390 0.280 2.600 0.730 ;
        RECT 3.230 0.280 3.480 0.730 ;
        RECT 4.110 0.280 4.360 0.730 ;
        RECT 4.990 0.280 5.240 0.730 ;
        RECT 5.870 0.280 6.120 0.730 ;
        RECT 6.760 0.700 7.200 0.730 ;
        RECT 6.760 0.280 7.010 0.700 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.570 1.680 0.830 2.460 ;
        RECT 1.440 1.680 1.710 2.460 ;
        RECT 0.570 1.510 2.220 1.680 ;
        RECT 2.050 1.340 2.220 1.510 ;
        RECT 2.050 1.070 6.520 1.340 ;
        RECT 2.050 0.900 2.220 1.070 ;
        RECT 0.570 0.720 2.220 0.900 ;
        RECT 0.570 0.280 0.820 0.720 ;
        RECT 1.450 0.280 1.700 0.720 ;
  END
END sky130_as_sc_hs__clkbuff_11

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_3
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.110 -0.075 0.380 0.220 ;
        RECT 0.110 -0.110 0.360 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.980 0.580 1.580 ;
        RECT 0.140 0.105 1.210 0.980 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.140 1.830 1.210 2.630 ;
        RECT 0.830 1.150 1.170 1.830 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
END sky130_as_sc_hs__decap_3

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.110 0.240 1.730 1.020 ;
        RECT 0.130 0.220 1.600 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.170 1.850 1.670 2.630 ;
        RECT 1.270 1.180 1.610 1.850 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.240 0.900 0.580 1.580 ;
        RECT 0.180 0.105 1.660 0.900 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_4

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__decap_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__decap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.220 7.120 1.020 ;
        RECT 0.120 -0.110 0.520 0.220 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
        RECT 0.360 1.690 6.980 2.630 ;
        RECT 0.600 1.340 0.850 1.690 ;
        RECT 0.560 1.140 0.890 1.340 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 6.390 0.940 6.720 1.520 ;
        RECT 0.360 0.105 6.970 0.940 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__decap_16

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.240 8.710 1.020 ;
        RECT 0.110 0.220 8.040 0.240 ;
        RECT 0.110 -0.075 0.410 0.220 ;
        RECT 0.110 -0.100 0.320 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 8.740 2.810 ;
        RECT 0.620 2.090 0.790 2.630 ;
        RECT 1.610 2.070 1.780 2.630 ;
        RECT 3.990 2.080 4.160 2.630 ;
        RECT 6.510 2.080 6.680 2.630 ;
        RECT 7.485 1.860 7.655 2.630 ;
        RECT 8.345 1.860 8.515 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.620 0.105 0.790 0.640 ;
        RECT 1.610 0.105 1.780 0.750 ;
        RECT 4.030 0.105 4.200 0.650 ;
        RECT 6.520 0.105 6.690 0.650 ;
        RECT 7.485 0.105 7.655 0.840 ;
        RECT 8.345 0.105 8.515 0.840 ;
        RECT 0.000 -0.085 8.740 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.169500 ;
    PORT
      LAYER li1 ;
        RECT 0.120 1.220 0.440 1.580 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.350000 ;
    PORT
      LAYER li1 ;
        RECT 7.890 1.690 8.110 2.420 ;
        RECT 7.690 1.150 8.110 1.690 ;
        RECT 7.890 0.300 8.110 1.150 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 1.580 0.920 1.910 1.680 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.190 1.920 0.360 2.440 ;
        RECT 1.060 1.920 1.230 2.440 ;
        RECT 0.190 1.750 0.780 1.920 ;
        RECT 1.060 1.750 1.410 1.920 ;
        RECT 0.610 1.450 0.780 1.750 ;
        RECT 1.210 1.590 1.410 1.750 ;
        RECT 0.610 1.180 1.070 1.450 ;
        RECT 0.610 0.980 0.780 1.180 ;
        RECT 1.240 1.010 1.410 1.590 ;
        RECT 0.190 0.810 0.780 0.980 ;
        RECT 1.060 0.840 1.410 1.010 ;
        RECT 0.190 0.280 0.360 0.810 ;
        RECT 1.060 0.280 1.230 0.840 ;
        RECT 2.080 0.280 2.250 2.450 ;
        RECT 2.550 2.210 2.970 2.380 ;
        RECT 2.420 1.560 2.630 1.890 ;
        RECT 2.800 1.780 2.970 2.210 ;
        RECT 4.170 1.780 4.380 1.850 ;
        RECT 2.800 1.610 4.380 1.780 ;
        RECT 2.420 1.050 2.630 1.380 ;
        RECT 2.800 0.880 2.970 1.610 ;
        RECT 4.170 1.520 4.380 1.610 ;
        RECT 3.800 1.230 4.010 1.310 ;
        RECT 4.550 1.230 4.720 2.450 ;
        RECT 5.030 2.210 5.450 2.380 ;
        RECT 4.890 1.560 5.100 1.890 ;
        RECT 5.280 1.790 5.450 2.210 ;
        RECT 6.940 2.030 7.200 2.460 ;
        RECT 6.670 1.790 6.860 1.850 ;
        RECT 5.280 1.620 6.860 1.790 ;
        RECT 2.710 0.710 2.970 0.880 ;
        RECT 3.300 0.830 3.510 1.160 ;
        RECT 3.800 1.060 4.720 1.230 ;
        RECT 3.800 0.980 4.010 1.060 ;
        RECT 2.710 0.600 2.880 0.710 ;
        RECT 2.550 0.430 2.880 0.600 ;
        RECT 4.550 0.290 4.720 1.060 ;
        RECT 4.900 1.050 5.110 1.380 ;
        RECT 5.280 0.880 5.450 1.620 ;
        RECT 6.670 1.520 6.860 1.620 ;
        RECT 7.030 1.590 7.200 2.030 ;
        RECT 6.280 1.230 6.490 1.310 ;
        RECT 7.030 1.260 7.470 1.590 ;
        RECT 7.030 1.230 7.200 1.260 ;
        RECT 5.190 0.710 5.450 0.880 ;
        RECT 5.790 0.830 6.000 1.160 ;
        RECT 6.280 1.060 7.200 1.230 ;
        RECT 6.280 0.980 6.490 1.060 ;
        RECT 7.030 0.790 7.200 1.060 ;
        RECT 5.190 0.600 5.360 0.710 ;
        RECT 5.030 0.430 5.360 0.600 ;
        RECT 6.955 0.670 7.200 0.790 ;
        RECT 6.955 0.280 7.160 0.670 ;
      LAYER met1 ;
        RECT 1.170 1.610 4.390 1.840 ;
        RECT 4.840 1.610 5.990 1.840 ;
        RECT 1.170 1.590 1.470 1.610 ;
        RECT 0.760 1.180 1.070 1.450 ;
        RECT 0.760 0.630 0.900 1.180 ;
        RECT 2.380 1.100 2.690 1.340 ;
        RECT 3.300 1.190 3.520 1.610 ;
        RECT 4.210 1.320 4.390 1.610 ;
        RECT 4.970 1.330 5.110 1.340 ;
        RECT 4.860 1.320 5.170 1.330 ;
        RECT 2.500 1.090 2.690 1.100 ;
        RECT 2.500 0.640 2.640 1.090 ;
        RECT 3.290 0.820 3.540 1.190 ;
        RECT 4.210 1.150 5.170 1.320 ;
        RECT 5.770 1.190 5.990 1.610 ;
        RECT 4.860 1.090 5.170 1.150 ;
        RECT 4.970 1.050 5.110 1.090 ;
        RECT 5.760 0.820 6.030 1.190 ;
        RECT 5.860 0.640 6.000 0.820 ;
        RECT 2.470 0.630 6.000 0.640 ;
        RECT 0.760 0.490 6.000 0.630 ;
  END
END sky130_as_sc_hs__dfxtp_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__diode_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.220 0.870 1.020 ;
        RECT 0.210 -0.075 0.390 0.220 ;
    END
  END VNB
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.441000 ;
    PORT
      LAYER li1 ;
        RECT 0.190 0.290 0.740 2.450 ;
    END
  END DIODE
END sky130_as_sc_hs__diode_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 0.920 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__fill_4

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_as_sc_hs__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.210 0.360 0.450 2.360 ;
  END
END sky130_as_sc_hs__fill_8

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__fill_16
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 7.360 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 7.360 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.730 2.020 0.970 2.260 ;
        RECT 0.490 1.780 1.210 2.020 ;
        RECT 0.490 1.300 0.730 1.780 ;
        RECT 0.970 1.300 1.210 1.780 ;
        RECT 1.690 1.540 1.930 2.260 ;
        RECT 3.130 1.540 3.370 2.260 ;
        RECT 4.090 2.020 4.330 2.260 ;
        RECT 1.690 1.300 2.170 1.540 ;
        RECT 0.490 1.060 1.210 1.300 ;
        RECT 0.250 0.820 0.730 1.060 ;
        RECT 0.970 0.820 1.450 1.060 ;
        RECT 0.250 0.340 0.490 0.820 ;
        RECT 1.210 0.340 1.450 0.820 ;
        RECT 1.930 0.820 2.170 1.300 ;
        RECT 2.410 0.820 2.650 1.540 ;
        RECT 2.890 1.300 3.370 1.540 ;
        RECT 3.850 1.780 4.570 2.020 ;
        RECT 3.850 1.300 4.090 1.780 ;
        RECT 4.330 1.300 4.570 1.780 ;
        RECT 5.050 1.540 5.290 2.260 ;
        RECT 6.490 1.540 6.730 2.260 ;
        RECT 5.050 1.300 5.530 1.540 ;
        RECT 2.890 0.820 3.130 1.300 ;
        RECT 3.850 1.060 4.570 1.300 ;
        RECT 1.930 0.580 3.130 0.820 ;
        RECT 3.610 0.820 4.090 1.060 ;
        RECT 4.330 0.820 4.810 1.060 ;
        RECT 2.170 0.340 2.410 0.580 ;
        RECT 2.650 0.340 2.890 0.580 ;
        RECT 3.610 0.340 3.850 0.820 ;
        RECT 4.570 0.340 4.810 0.820 ;
        RECT 5.290 0.820 5.530 1.300 ;
        RECT 5.770 0.820 6.010 1.540 ;
        RECT 6.250 1.300 6.730 1.540 ;
        RECT 6.250 0.820 6.490 1.300 ;
        RECT 5.290 0.580 6.490 0.820 ;
        RECT 5.530 0.340 5.770 0.580 ;
        RECT 6.010 0.340 6.250 0.580 ;
  END
END sky130_as_sc_hs__fill_16

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.220 1.600 1.020 ;
        RECT 0.120 -0.075 0.380 0.220 ;
        RECT 0.120 -0.110 0.350 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.840 2.810 ;
        RECT 0.320 1.490 0.570 2.630 ;
        RECT 1.320 1.490 1.570 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.310 0.105 0.560 0.880 ;
        RECT 1.310 0.105 1.530 0.870 ;
        RECT 0.000 -0.085 1.840 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490500 ;
    PORT
      LAYER li1 ;
        RECT 0.820 0.310 1.070 2.430 ;
    END
  END Y
  PIN A
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.654000 ;
    PORT
      LAYER li1 ;
        RECT 0.320 1.050 0.650 1.320 ;
    END
  END A
END sky130_as_sc_hs__inv_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__inv_4
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.890 2.710 1.020 ;
        RECT 0.120 0.240 2.760 0.890 ;
        RECT 0.120 0.220 2.710 0.240 ;
        RECT 0.120 -0.075 0.380 0.220 ;
        RECT 1.480 0.110 2.230 0.220 ;
        RECT 2.050 -0.075 2.230 0.110 ;
        RECT 0.120 -0.110 0.350 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.760 2.810 ;
        RECT 0.320 1.620 0.570 2.630 ;
        RECT 1.320 1.490 1.570 2.630 ;
        RECT 2.320 1.490 2.530 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.310 0.105 0.560 0.780 ;
        RECT 1.310 0.105 1.530 0.870 ;
        RECT 2.310 0.105 2.520 0.890 ;
        RECT 0.000 -0.085 2.760 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.981000 ;
    PORT
      LAYER li1 ;
        RECT 0.820 1.320 1.070 2.430 ;
        RECT 1.780 1.320 2.030 2.430 ;
        RECT 0.820 1.120 2.030 1.320 ;
        RECT 0.820 0.310 1.070 1.120 ;
        RECT 1.780 0.310 2.030 1.120 ;
    END
  END Y
  PIN A
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.308000 ;
    PORT
      LAYER li1 ;
        RECT 0.320 0.950 0.650 1.450 ;
    END
  END A
END sky130_as_sc_hs__inv_4

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__mux2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.110 0.240 4.100 1.020 ;
        RECT 0.130 0.220 1.600 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 4.330 2.910 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 4.140 2.810 ;
        RECT 0.605 2.180 0.775 2.630 ;
        RECT 2.870 1.940 3.130 2.630 ;
        RECT 3.815 1.860 3.985 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.105 0.775 0.590 ;
        RECT 2.760 0.105 3.140 0.540 ;
        RECT 3.815 0.105 3.985 0.940 ;
        RECT 0.000 -0.085 4.140 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 2.080 1.750 2.350 1.810 ;
        RECT 1.740 1.480 2.350 1.750 ;
        RECT 0.450 1.130 0.680 1.140 ;
        RECT 0.450 1.120 1.490 1.130 ;
        RECT 1.740 1.120 1.920 1.480 ;
        RECT 0.450 0.950 1.920 1.120 ;
        RECT 0.450 0.810 1.490 0.950 ;
        RECT 1.240 0.800 1.490 0.810 ;
    END
  END S
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156750 ;
    PORT
      LAYER li1 ;
        RECT 0.670 1.340 1.000 1.670 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.165750 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.050 2.690 1.310 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.410200 ;
    PORT
      LAYER li1 ;
        RECT 3.385 1.690 3.555 2.430 ;
        RECT 3.385 1.120 3.830 1.690 ;
        RECT 3.385 0.280 3.555 1.120 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 2.010 0.345 2.440 ;
        RECT 1.570 2.150 1.990 2.380 ;
        RECT 1.570 2.080 2.700 2.150 ;
        RECT 0.175 1.840 1.410 2.010 ;
        RECT 1.630 1.980 2.700 2.080 ;
        RECT 0.175 1.530 0.345 1.840 ;
        RECT 0.110 1.340 0.345 1.530 ;
        RECT 1.240 1.720 1.410 1.840 ;
        RECT 2.530 1.730 2.700 1.980 ;
        RECT 1.240 1.390 1.510 1.720 ;
        RECT 2.530 1.560 3.150 1.730 ;
        RECT 2.860 1.540 3.150 1.560 ;
        RECT 0.110 0.660 0.280 1.340 ;
        RECT 2.860 1.210 3.210 1.540 ;
        RECT 2.860 0.880 3.030 1.210 ;
        RECT 2.410 0.710 3.030 0.880 ;
        RECT 0.110 0.500 0.345 0.660 ;
        RECT 2.410 0.620 2.590 0.710 ;
        RECT 0.175 0.290 0.345 0.500 ;
        RECT 1.480 0.450 2.590 0.620 ;
        RECT 1.480 0.290 1.920 0.450 ;
  END
END sky130_as_sc_hs__mux2_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.880 3.630 1.020 ;
        RECT 0.000 0.240 3.630 0.880 ;
        RECT 0.010 0.220 1.370 0.240 ;
        RECT 1.490 0.230 3.630 0.240 ;
        RECT 1.510 0.220 2.980 0.230 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
        RECT 1.510 -0.100 1.830 0.220 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.300 0.105 0.540 0.830 ;
        RECT 1.940 0.105 2.200 0.540 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.300 1.650 0.540 2.630 ;
        RECT 1.280 1.600 1.520 2.630 ;
        RECT 2.190 1.920 2.600 2.630 ;
        RECT 3.250 1.920 3.480 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    PORT
      LAYER li1 ;
        RECT 3.280 1.370 3.460 1.750 ;
        RECT 3.150 1.040 3.460 1.370 ;
        RECT 3.280 0.840 3.460 1.040 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699800 ;
    PORT
      LAYER li1 ;
        RECT 1.720 1.750 1.960 2.430 ;
        RECT 2.810 1.750 3.050 2.430 ;
        RECT 1.720 1.530 3.050 1.750 ;
        RECT 2.370 1.270 2.610 1.530 ;
        RECT 2.370 1.050 2.980 1.270 ;
        RECT 2.760 0.870 2.980 1.050 ;
        RECT 2.760 0.620 3.100 0.870 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.250 1.060 0.600 1.400 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.770 1.340 1.000 2.460 ;
        RECT 0.770 1.050 2.200 1.340 ;
        RECT 0.770 0.290 1.000 1.050 ;
        RECT 1.530 0.710 2.590 0.880 ;
        RECT 1.530 0.280 1.760 0.710 ;
        RECT 2.380 0.450 2.590 0.710 ;
        RECT 3.250 0.450 3.580 0.540 ;
        RECT 2.380 0.280 3.580 0.450 ;
  END
END sky130_as_sc_hs__nand2b_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__and2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.240 2.250 1.020 ;
        RECT 0.130 0.220 1.600 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 0.175 1.600 0.345 2.630 ;
        RECT 1.035 1.950 1.205 2.630 ;
        RECT 1.870 2.250 2.210 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.035 0.105 1.205 0.880 ;
        RECT 1.955 0.105 2.125 0.600 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.090 0.370 1.430 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.070 1.105 1.410 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.456750 ;
    PORT
      LAYER li1 ;
        RECT 1.515 2.080 1.685 2.450 ;
        RECT 1.515 1.950 2.000 2.080 ;
        RECT 1.560 1.910 2.000 1.950 ;
        RECT 1.700 0.920 2.000 1.910 ;
        RECT 1.515 0.770 2.000 0.920 ;
        RECT 1.515 0.750 1.870 0.770 ;
        RECT 1.515 0.280 1.685 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.605 1.810 0.775 2.460 ;
        RECT 0.540 1.780 0.775 1.810 ;
        RECT 0.540 1.600 1.445 1.780 ;
        RECT 0.540 0.920 0.710 1.600 ;
        RECT 1.275 1.440 1.445 1.600 ;
        RECT 1.275 1.090 1.530 1.440 ;
        RECT 0.170 0.750 0.710 0.920 ;
        RECT 0.175 0.280 0.345 0.750 ;
  END
END sky130_as_sc_hs__and2_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nand3_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.240 3.670 1.020 ;
        RECT 0.110 0.230 2.250 0.240 ;
        RECT 0.130 0.220 1.600 0.230 ;
        RECT 2.310 0.220 3.670 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
        RECT 2.430 -0.075 2.680 0.220 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.175 1.590 0.345 2.630 ;
        RECT 1.035 1.920 1.205 2.630 ;
        RECT 1.900 1.920 2.610 2.630 ;
        RECT 3.325 1.920 3.495 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.560 0.105 0.820 0.540 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.050 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.610 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.060 2.630 1.340 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.942200 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.750 0.800 2.410 ;
        RECT 1.430 1.750 1.670 2.430 ;
        RECT 2.860 1.750 3.100 2.430 ;
        RECT 0.580 1.530 3.100 1.750 ;
        RECT 2.810 0.890 3.100 1.530 ;
        RECT 2.810 0.620 3.150 0.890 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.150 0.710 1.210 0.880 ;
        RECT 0.150 0.280 0.380 0.710 ;
        RECT 1.000 0.450 1.210 0.710 ;
        RECT 1.380 0.680 2.630 0.890 ;
        RECT 1.380 0.620 1.720 0.680 ;
        RECT 1.850 0.450 2.180 0.510 ;
        RECT 1.000 0.280 2.180 0.450 ;
        RECT 2.420 0.450 2.630 0.680 ;
        RECT 3.315 0.450 3.580 0.570 ;
        RECT 2.420 0.280 3.580 0.450 ;
  END
END sky130_as_sc_hs__nand3_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.240 2.250 1.020 ;
        RECT 0.110 0.230 2.250 0.240 ;
        RECT 0.130 0.220 1.600 0.230 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 0.550 1.970 0.830 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.860 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.900 0.105 2.070 0.540 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.060 0.980 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER li1 ;
        RECT 1.190 1.060 1.610 1.340 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.610400 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.750 1.680 2.070 ;
        RECT 1.420 1.520 2.160 1.750 ;
        RECT 1.780 0.890 2.160 1.520 ;
        RECT 0.570 0.710 2.160 0.890 ;
        RECT 0.570 0.280 0.790 0.710 ;
        RECT 1.440 0.280 1.660 0.710 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.150 1.800 0.380 2.460 ;
        RECT 1.000 2.240 2.160 2.460 ;
        RECT 1.000 1.800 1.240 2.240 ;
        RECT 1.910 1.920 2.160 2.240 ;
        RECT 0.150 1.570 1.240 1.800 ;
  END
END sky130_as_sc_hs__nor2_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.240 3.670 1.020 ;
        RECT 0.110 0.230 3.670 0.240 ;
        RECT 0.130 0.220 1.600 0.230 ;
        RECT 2.310 0.220 3.670 0.230 ;
        RECT 0.130 -0.100 0.450 0.220 ;
        RECT 2.430 -0.075 2.680 0.220 ;
        RECT 2.430 -0.100 2.630 -0.075 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 3.680 2.810 ;
        RECT 0.550 1.970 0.830 2.630 ;
        RECT 3.270 1.590 3.460 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.490 3.680 2.960 ;
        RECT 0.000 2.480 2.370 2.490 ;
        RECT 2.770 2.480 3.680 2.490 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.860 ;
        RECT 1.035 0.105 1.205 0.540 ;
        RECT 1.900 0.105 2.070 0.830 ;
        RECT 3.280 0.105 3.450 0.850 ;
        RECT 0.000 -0.085 3.680 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 3.870 2.910 ;
    END
  END VPB
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.442500 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.060 0.980 1.340 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.590800 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.400 1.680 2.070 ;
        RECT 1.150 1.210 1.680 1.400 ;
        RECT 1.150 0.890 1.380 1.210 ;
        RECT 0.570 0.710 1.660 0.890 ;
        RECT 0.570 0.280 0.790 0.710 ;
        RECT 1.440 0.280 1.660 0.710 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225750 ;
    PORT
      LAYER li1 ;
        RECT 3.230 1.020 3.530 1.420 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 0.150 1.800 0.380 2.460 ;
        RECT 1.000 2.240 2.130 2.460 ;
        RECT 1.000 1.800 1.240 2.240 ;
        RECT 1.850 1.920 2.130 2.240 ;
        RECT 0.150 1.570 1.240 1.800 ;
        RECT 1.870 1.240 2.080 1.360 ;
        RECT 2.810 1.240 3.060 2.430 ;
        RECT 1.870 1.020 3.060 1.240 ;
        RECT 1.870 1.000 2.080 1.020 ;
        RECT 2.810 0.310 3.060 1.020 ;
  END
END sky130_as_sc_hs__nor2b_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__or2_2
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.240 2.250 1.020 ;
        RECT 0.130 0.220 1.600 0.240 ;
        RECT 0.130 -0.100 0.450 0.220 ;
    END
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.490 2.910 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 2.300 2.810 ;
        RECT 1.035 1.950 1.205 2.630 ;
        RECT 1.870 2.250 2.210 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.105 0.345 0.920 ;
        RECT 1.035 0.105 1.205 0.860 ;
        RECT 1.955 0.105 2.125 0.600 ;
        RECT 0.000 -0.085 2.300 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.090 0.370 1.430 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.236250 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.030 1.105 1.440 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.456750 ;
    PORT
      LAYER li1 ;
        RECT 1.515 2.080 1.685 2.450 ;
        RECT 1.515 1.950 2.000 2.080 ;
        RECT 1.560 1.910 2.000 1.950 ;
        RECT 1.700 0.920 2.000 1.910 ;
        RECT 1.515 0.770 2.000 0.920 ;
        RECT 1.515 0.750 1.870 0.770 ;
        RECT 1.515 0.280 1.685 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.175 1.780 0.345 2.460 ;
        RECT 0.175 1.610 1.445 1.780 ;
        RECT 0.175 1.600 0.710 1.610 ;
        RECT 0.540 0.860 0.710 1.600 ;
        RECT 1.275 1.440 1.445 1.610 ;
        RECT 1.275 1.090 1.530 1.440 ;
        RECT 0.540 0.280 0.775 0.860 ;
  END
END sky130_as_sc_hs__or2_2

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tap_1
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.000 2.630 0.460 2.810 ;
        RECT 0.110 1.460 0.340 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.220 0.430 1.020 ;
        RECT 0.090 -0.120 0.400 0.220 ;
      LAYER li1 ;
        RECT 0.120 0.105 0.340 1.000 ;
        RECT 0.000 -0.085 0.460 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
END sky130_as_sc_hs__tap_1

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tieh
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.730 1.840 1.040 2.630 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 0.380 1.040 1.630 ;
    END
  END ONE
END sky130_as_sc_hs__tieh

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_as_sc_hs__tiel
  CLASS CORE ;
  FOREIGN sky130_as_sc_hs__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.220 1.370 1.020 ;
        RECT 0.130 -0.075 0.380 0.220 ;
        RECT 0.130 -0.100 0.330 -0.075 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 1.570 2.910 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.105 1.040 0.860 ;
        RECT 0.000 -0.085 1.380 0.105 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN ZERO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.300 1.140 1.040 2.390 ;
    END
  END ZERO
END sky130_as_sc_hs__tiel
END LIBRARY
