magic
tech sky130A
magscale 1 2
timestamp 1738764062
<< nwell >>
rect -38 262 866 582
<< pwell >>
rect 0 26 828 204
rect 22 -20 90 26
<< pmos >>
rect 80 323 110 496
rect 168 323 198 496
rect 256 323 286 496
rect 344 323 374 496
rect 432 323 462 496
rect 519 323 549 496
rect 605 323 635 496
rect 691 323 721 496
<< nmoslvt >>
rect 80 49 110 179
rect 168 49 198 179
rect 256 49 286 179
rect 344 49 374 179
rect 432 49 462 179
rect 519 49 549 179
rect 605 49 635 179
rect 691 49 721 179
<< ndiff >>
rect 27 140 80 179
rect 27 76 35 140
rect 69 76 80 140
rect 27 49 80 76
rect 110 170 168 179
rect 110 72 121 170
rect 155 72 168 170
rect 110 49 168 72
rect 198 171 256 179
rect 198 58 209 171
rect 243 58 256 171
rect 198 49 256 58
rect 286 171 344 179
rect 286 72 298 171
rect 332 72 344 171
rect 286 49 344 72
rect 374 120 432 179
rect 374 72 386 120
rect 420 72 432 120
rect 374 49 432 72
rect 462 171 519 179
rect 462 72 474 171
rect 508 72 519 171
rect 462 49 519 72
rect 549 166 605 179
rect 549 57 560 166
rect 594 57 605 166
rect 549 49 605 57
rect 635 171 691 179
rect 635 72 646 171
rect 680 72 691 171
rect 635 49 691 72
rect 721 170 801 179
rect 721 57 736 170
rect 770 57 801 170
rect 721 49 801 57
<< pdiff >>
rect 27 484 80 496
rect 27 350 35 484
rect 69 350 80 484
rect 27 323 80 350
rect 110 476 168 496
rect 110 331 121 476
rect 155 331 168 476
rect 110 323 168 331
rect 198 488 256 496
rect 198 346 209 488
rect 243 346 256 488
rect 198 323 256 346
rect 286 476 344 496
rect 286 354 298 476
rect 332 354 344 476
rect 286 323 344 354
rect 374 474 432 496
rect 374 406 386 474
rect 420 406 432 474
rect 374 323 432 406
rect 462 474 519 496
rect 462 354 474 474
rect 508 354 519 474
rect 462 323 519 354
rect 549 488 605 496
rect 549 342 560 488
rect 594 342 605 488
rect 549 323 605 342
rect 635 474 691 496
rect 635 331 646 474
rect 680 331 691 474
rect 635 323 691 331
rect 721 488 801 496
rect 721 342 734 488
rect 768 342 801 488
rect 721 323 801 342
<< ndiffc >>
rect 35 76 69 140
rect 121 72 155 170
rect 209 58 243 171
rect 298 72 332 171
rect 386 72 420 120
rect 474 72 508 171
rect 560 57 594 166
rect 646 72 680 171
rect 736 57 770 170
<< pdiffc >>
rect 35 350 69 484
rect 121 331 155 476
rect 209 346 243 488
rect 298 354 332 476
rect 386 406 420 474
rect 474 354 508 474
rect 560 342 594 488
rect 646 331 680 474
rect 734 342 768 488
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 519 496 549 522
rect 605 496 635 522
rect 691 496 721 522
rect 80 296 110 323
rect 168 296 198 323
rect 256 300 286 323
rect 28 276 198 296
rect 28 242 44 276
rect 78 242 198 276
rect 28 226 198 242
rect 240 292 296 300
rect 344 292 374 323
rect 432 292 462 323
rect 519 292 549 323
rect 605 292 635 323
rect 691 292 721 323
rect 240 276 721 292
rect 240 242 250 276
rect 284 242 721 276
rect 240 226 296 242
rect 80 179 110 226
rect 168 179 198 226
rect 256 179 286 226
rect 344 179 374 242
rect 432 179 462 242
rect 519 179 549 242
rect 605 179 635 242
rect 691 179 721 242
rect 80 23 110 49
rect 168 23 198 49
rect 256 23 286 49
rect 344 23 374 49
rect 432 23 462 49
rect 519 23 549 49
rect 605 23 635 49
rect 691 23 721 49
<< polycont >>
rect 44 242 78 276
rect 250 242 284 276
<< locali >>
rect 0 561 828 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 526 828 527
rect 35 484 69 526
rect 35 334 69 350
rect 120 476 156 492
rect 120 331 121 476
rect 155 331 156 476
rect 31 276 84 296
rect 31 242 44 276
rect 78 242 84 276
rect 31 226 84 242
rect 120 284 156 331
rect 209 488 243 526
rect 209 330 243 346
rect 298 476 332 492
rect 386 474 420 526
rect 386 390 420 406
rect 474 474 508 490
rect 332 354 356 372
rect 298 338 356 354
rect 322 304 356 338
rect 474 304 508 354
rect 560 488 594 526
rect 560 326 594 342
rect 646 474 680 490
rect 238 284 284 296
rect 120 276 284 284
rect 120 244 250 276
rect 120 170 156 244
rect 238 242 250 244
rect 238 226 284 242
rect 322 292 508 304
rect 646 292 680 331
rect 734 488 768 526
rect 734 326 768 342
rect 322 226 680 292
rect 35 140 69 158
rect 35 21 69 76
rect 120 72 121 170
rect 155 72 156 170
rect 120 56 156 72
rect 209 171 243 192
rect 322 188 356 226
rect 209 21 243 58
rect 298 171 356 188
rect 332 154 356 171
rect 474 171 508 226
rect 298 56 332 72
rect 386 120 420 136
rect 386 21 420 72
rect 474 56 508 72
rect 560 166 594 182
rect 560 21 594 57
rect 646 171 680 226
rect 646 56 680 72
rect 736 170 770 190
rect 736 21 770 57
rect 0 17 828 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_6
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali 357 255 391 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 374 272 374 272 0 FreeSans 200 0 0 0 Y
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_6.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 828 216
string MASKHINTS_NSDM 0 -38 828 204
string MASKHINTS_PSDM 0 272 828 582
<< end >>
