magic
tech sky130A
magscale 1 2
timestamp 1739628591
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 10 48 450 204
rect 26 44 320 48
rect 26 26 90 44
rect 26 22 110 26
rect 26 -20 90 22
<< pmos >>
rect 80 314 110 496
rect 166 314 196 496
rect 262 314 292 496
rect 350 314 380 496
<< nmoslvt >>
rect 80 48 110 184
rect 166 48 196 184
rect 262 48 292 184
rect 350 48 380 184
<< ndiff >>
rect 27 166 80 184
rect 27 72 35 166
rect 69 72 80 166
rect 27 48 80 72
rect 110 48 166 184
rect 196 156 262 184
rect 196 72 207 156
rect 241 72 262 156
rect 196 48 262 72
rect 292 166 350 184
rect 292 72 303 166
rect 337 72 350 166
rect 292 48 350 72
rect 380 102 433 184
rect 380 61 391 102
rect 425 61 433 102
rect 380 48 433 61
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 314 80 336
rect 110 476 166 496
rect 110 348 121 476
rect 155 348 166 476
rect 110 314 166 348
rect 196 488 262 496
rect 196 406 207 488
rect 241 406 262 488
rect 196 314 262 406
rect 292 474 350 496
rect 292 406 303 474
rect 337 406 350 474
rect 292 314 350 406
rect 380 484 433 496
rect 380 450 391 484
rect 425 450 433 484
rect 380 314 433 450
<< ndiffc >>
rect 35 72 69 166
rect 207 72 241 156
rect 303 72 337 166
rect 391 61 425 102
<< pdiffc >>
rect 35 336 69 476
rect 121 348 155 476
rect 207 406 241 488
rect 303 406 337 474
rect 391 450 425 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 262 496 292 522
rect 350 496 380 522
rect 80 284 110 314
rect 30 266 110 284
rect 30 232 40 266
rect 74 232 110 266
rect 30 216 110 232
rect 80 184 110 216
rect 166 284 196 314
rect 262 288 292 314
rect 350 288 380 314
rect 166 266 220 284
rect 166 232 176 266
rect 210 232 220 266
rect 166 212 220 232
rect 262 266 380 288
rect 262 232 272 266
rect 306 232 380 266
rect 262 216 380 232
rect 166 184 196 212
rect 262 184 292 216
rect 350 184 380 216
rect 80 22 110 48
rect 166 22 196 48
rect 262 22 292 48
rect 350 22 380 48
<< polycont >>
rect 40 232 74 266
rect 176 232 210 266
rect 272 232 306 266
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 35 476 69 526
rect 121 476 155 492
rect 35 320 69 336
rect 108 348 121 362
rect 207 488 241 526
rect 207 390 241 406
rect 303 474 337 490
rect 374 484 442 526
rect 374 450 391 484
rect 425 450 442 484
rect 337 406 400 416
rect 303 390 400 406
rect 312 382 400 390
rect 155 348 289 356
rect 108 320 289 348
rect 30 266 74 286
rect 30 232 40 266
rect 30 216 74 232
rect 108 182 142 320
rect 255 288 289 320
rect 176 266 221 282
rect 210 232 221 266
rect 176 214 221 232
rect 255 266 306 288
rect 255 232 272 266
rect 255 216 306 232
rect 340 182 400 382
rect 34 166 142 182
rect 34 148 35 166
rect 69 148 142 166
rect 207 156 241 176
rect 35 56 69 72
rect 207 21 241 72
rect 303 166 400 182
rect 337 154 400 166
rect 337 148 374 154
rect 303 56 337 72
rect 391 102 425 118
rect 391 21 425 61
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
flabel locali 187 221 221 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 204 238 204 238 0 FreeSans 200 0 0 0 B
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__and2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 220
string MASKHINTS_NSDM 0 -38 460 209
string MASKHINTS_PSDM 0 289 460 582
<< end >>
