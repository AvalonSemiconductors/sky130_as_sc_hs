magic
tech sky130A
magscale 1 2
timestamp 1738971918
<< nwell >>
rect -38 262 1050 582
<< pwell >>
rect 0 28 1012 204
rect 0 22 736 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 252 298 282 496
rect 338 298 368 496
rect 578 298 608 496
rect 664 298 694 496
rect 750 298 780 496
rect 836 298 866 496
<< nmoslvt >>
rect 80 49 110 178
rect 166 49 196 178
rect 252 49 282 178
rect 338 49 368 178
rect 578 49 608 178
rect 664 49 694 178
rect 750 49 780 178
rect 836 49 866 178
<< ndiff >>
rect 27 162 80 178
rect 27 62 35 162
rect 69 62 80 162
rect 27 49 80 62
rect 110 162 166 178
rect 110 72 121 162
rect 155 72 166 162
rect 110 49 166 72
rect 196 92 252 178
rect 196 58 207 92
rect 241 58 252 92
rect 196 49 252 58
rect 282 162 338 178
rect 282 72 293 162
rect 327 72 338 162
rect 282 49 338 72
rect 368 92 426 178
rect 368 58 379 92
rect 413 58 426 92
rect 368 49 426 58
rect 480 170 578 178
rect 480 136 533 170
rect 567 136 578 170
rect 480 49 578 136
rect 608 94 664 178
rect 608 60 619 94
rect 653 60 664 94
rect 608 49 664 60
rect 694 162 750 178
rect 694 76 705 162
rect 739 76 750 162
rect 694 49 750 76
rect 780 170 836 178
rect 780 136 791 170
rect 825 136 836 170
rect 780 49 836 136
rect 866 162 960 178
rect 866 76 884 162
rect 918 76 960 162
rect 866 49 960 76
<< pdiff >>
rect 27 476 80 496
rect 27 320 35 476
rect 69 320 80 476
rect 27 298 80 320
rect 110 488 166 496
rect 110 388 121 488
rect 155 388 166 488
rect 110 298 166 388
rect 196 476 252 496
rect 196 320 207 476
rect 241 320 252 476
rect 196 298 252 320
rect 282 406 338 496
rect 282 318 293 406
rect 327 318 338 406
rect 282 298 338 318
rect 368 468 426 496
rect 368 386 379 468
rect 413 386 426 468
rect 368 298 426 386
rect 480 488 578 496
rect 480 386 510 488
rect 544 386 578 488
rect 480 298 578 386
rect 608 476 664 496
rect 608 306 619 476
rect 653 306 664 476
rect 608 298 664 306
rect 694 488 750 496
rect 694 386 705 488
rect 739 386 750 488
rect 694 298 750 386
rect 780 474 836 496
rect 780 306 791 474
rect 825 306 836 474
rect 780 298 836 306
rect 866 488 960 496
rect 866 310 892 488
rect 926 310 960 488
rect 866 298 960 310
<< ndiffc >>
rect 35 62 69 162
rect 121 72 155 162
rect 207 58 241 92
rect 293 72 327 162
rect 379 58 413 92
rect 533 136 567 170
rect 619 60 653 94
rect 705 76 739 162
rect 791 136 825 170
rect 884 76 918 162
<< pdiffc >>
rect 35 320 69 476
rect 121 388 155 488
rect 207 320 241 476
rect 293 318 327 406
rect 379 386 413 468
rect 510 386 544 488
rect 619 306 653 476
rect 705 386 739 488
rect 791 306 825 474
rect 892 310 926 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 252 496 282 522
rect 338 496 368 522
rect 578 496 608 522
rect 664 496 694 522
rect 750 496 780 522
rect 836 496 866 522
rect 80 260 110 298
rect 166 260 196 298
rect 80 256 196 260
rect 78 250 196 256
rect 78 216 92 250
rect 126 216 196 250
rect 78 212 196 216
rect 80 204 196 212
rect 80 178 110 204
rect 166 178 196 204
rect 252 260 282 298
rect 338 260 368 298
rect 252 250 368 260
rect 252 216 268 250
rect 302 216 368 250
rect 252 204 368 216
rect 252 178 282 204
rect 338 178 368 204
rect 578 260 608 298
rect 664 260 694 298
rect 578 250 694 260
rect 578 216 594 250
rect 628 216 694 250
rect 578 204 694 216
rect 578 178 608 204
rect 664 178 694 204
rect 750 260 780 298
rect 836 260 866 298
rect 750 250 926 260
rect 750 216 876 250
rect 910 216 926 250
rect 750 204 926 216
rect 750 178 780 204
rect 836 178 866 204
rect 80 23 110 49
rect 166 23 196 49
rect 252 23 282 49
rect 338 23 368 49
rect 578 23 608 49
rect 664 23 694 49
rect 750 23 780 49
rect 836 23 866 49
<< polycont >>
rect 92 216 126 250
rect 268 216 302 250
rect 594 216 628 250
rect 876 216 910 250
<< locali >>
rect 0 561 1012 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 526 1012 527
rect 35 476 69 492
rect 121 488 155 526
rect 121 372 155 388
rect 207 476 413 492
rect 69 320 207 338
rect 241 468 413 476
rect 241 456 379 468
rect 35 304 241 320
rect 293 406 327 422
rect 379 370 413 386
rect 510 488 544 526
rect 510 370 544 386
rect 619 476 653 492
rect 327 318 619 336
rect 293 306 619 318
rect 705 488 739 526
rect 705 370 739 386
rect 774 474 825 490
rect 774 336 791 474
rect 653 306 791 336
rect 293 302 825 306
rect 76 250 142 256
rect 76 216 92 250
rect 126 216 142 250
rect 76 212 142 216
rect 252 250 318 256
rect 252 216 268 250
rect 302 216 318 250
rect 252 212 318 216
rect 578 250 644 256
rect 578 216 594 250
rect 628 216 644 250
rect 578 212 644 216
rect 35 162 69 178
rect 35 21 69 62
rect 121 162 482 178
rect 155 144 293 162
rect 121 56 155 72
rect 207 92 241 108
rect 207 21 241 58
rect 327 144 482 162
rect 293 56 327 72
rect 379 92 413 108
rect 448 96 482 144
rect 516 170 739 178
rect 516 136 533 170
rect 567 162 739 170
rect 567 144 705 162
rect 567 136 583 144
rect 619 96 653 110
rect 448 94 653 96
rect 448 62 619 94
rect 600 60 619 62
rect 653 60 670 94
rect 774 174 825 302
rect 892 488 926 526
rect 892 294 926 310
rect 860 250 926 256
rect 860 216 876 250
rect 910 216 926 250
rect 860 212 926 216
rect 774 170 842 174
rect 774 136 791 170
rect 825 136 842 170
rect 774 128 842 136
rect 884 162 918 178
rect 739 76 884 94
rect 705 60 918 76
rect 379 21 413 58
rect 0 17 1012 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ioa211_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1012 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 85 221 119 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali 102 238 102 238 0 FreeSans 200 0 0 0 A
flabel locali 272 221 306 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali 289 238 289 238 0 FreeSans 200 0 0 0 B
flabel locali 595 221 629 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali 612 238 612 238 0 FreeSans 200 0 0 0 C
flabel locali 884 221 918 255 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel locali 901 238 901 238 0 FreeSans 200 0 0 0 D
flabel locali 782 221 816 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali 799 238 799 238 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__ioa211_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1012 214
string MASKHINTS_NSDM 0 -38 1012 204
string MASKHINTS_PSDM 0 272 1012 582
<< end >>
