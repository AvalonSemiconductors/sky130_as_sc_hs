magic
tech sky130A
magscale 1 2
timestamp 1740281738
<< nwell >>
rect -38 262 498 582
<< pwell >>
rect 10 48 450 204
rect 26 44 320 48
rect 26 26 90 44
rect 26 22 110 26
rect 26 -20 90 22
<< pmos >>
rect 80 314 110 496
rect 166 314 196 496
rect 264 314 294 496
rect 350 314 380 496
<< nmoslvt >>
rect 80 48 110 184
rect 166 48 196 184
rect 264 48 294 184
rect 350 48 380 184
<< ndiff >>
rect 27 166 80 184
rect 27 72 35 166
rect 69 72 80 166
rect 27 48 80 72
rect 110 48 166 184
rect 196 156 264 184
rect 196 72 207 156
rect 241 72 264 156
rect 196 48 264 72
rect 294 166 350 184
rect 294 132 305 166
rect 339 132 350 166
rect 294 48 350 132
rect 380 102 433 184
rect 380 61 391 102
rect 425 61 433 102
rect 380 48 433 61
<< pdiff >>
rect 27 476 80 496
rect 27 336 35 476
rect 69 336 80 476
rect 27 314 80 336
rect 110 476 166 496
rect 110 348 121 476
rect 155 348 166 476
rect 110 314 166 348
rect 196 488 264 496
rect 196 406 207 488
rect 241 406 264 488
rect 196 314 264 406
rect 294 440 350 496
rect 294 406 305 440
rect 339 406 350 440
rect 294 314 350 406
rect 380 484 433 496
rect 380 450 391 484
rect 425 450 433 484
rect 380 314 433 450
<< ndiffc >>
rect 35 72 69 166
rect 207 72 241 156
rect 305 132 339 166
rect 391 61 425 102
<< pdiffc >>
rect 35 336 69 476
rect 121 348 155 476
rect 207 406 241 488
rect 305 406 339 440
rect 391 450 425 484
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 264 496 294 522
rect 350 496 380 522
rect 80 284 110 314
rect 30 266 110 284
rect 30 232 42 266
rect 76 232 110 266
rect 30 216 110 232
rect 80 184 110 216
rect 166 284 196 314
rect 264 288 294 314
rect 350 288 380 314
rect 166 266 222 284
rect 166 232 178 266
rect 212 232 222 266
rect 166 212 222 232
rect 264 266 380 288
rect 264 232 274 266
rect 308 232 380 266
rect 264 216 380 232
rect 166 184 196 212
rect 264 184 294 216
rect 350 184 380 216
rect 80 22 110 48
rect 166 22 196 48
rect 264 22 294 48
rect 350 22 380 48
<< polycont >>
rect 42 232 76 266
rect 178 232 212 266
rect 274 232 308 266
<< locali >>
rect 0 561 460 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 526 460 527
rect 35 476 69 526
rect 121 476 155 492
rect 35 320 69 336
rect 110 348 121 362
rect 207 488 241 526
rect 374 484 442 526
rect 207 390 241 406
rect 303 440 340 456
rect 374 450 391 484
rect 425 450 442 484
rect 303 406 305 440
rect 339 416 340 440
rect 339 406 392 416
rect 303 390 392 406
rect 312 382 392 390
rect 155 348 290 356
rect 110 320 290 348
rect 30 266 76 286
rect 30 232 42 266
rect 30 216 76 232
rect 110 182 144 320
rect 256 288 290 320
rect 178 266 222 282
rect 212 232 222 266
rect 178 214 222 232
rect 256 266 308 288
rect 256 232 274 266
rect 256 216 308 232
rect 342 182 392 382
rect 34 166 144 182
rect 34 148 35 166
rect 69 148 144 166
rect 207 156 241 176
rect 35 56 69 72
rect 303 166 392 182
rect 303 132 305 166
rect 339 154 392 166
rect 339 148 374 154
rect 303 116 339 132
rect 207 21 241 72
rect 391 102 425 118
rect 391 21 425 61
rect 0 17 460 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2_2
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 460 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 34 238 68 272 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel locali s 51 255 51 255 0 FreeSans 200 0 0 0 A
flabel locali s 357 221 391 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 238 375 238 0 FreeSans 200 0 0 0 Y
flabel locali s 357 340 391 374 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 375 357 375 357 0 FreeSans 200 0 0 0 Y
flabel locali 187 221 221 255 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel locali 204 238 204 238 0 FreeSans 200 0 0 0 B
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__and2_2.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 460 220
string MASKHINTS_NSDM 0 -38 460 209
string MASKHINTS_PSDM 0 289 460 582
<< end >>
