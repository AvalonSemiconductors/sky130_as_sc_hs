magic
tech sky130A
magscale 1 2
timestamp 1733757194
<< nwell >>
rect -38 262 130 582
<< locali >>
rect 0 561 92 562
rect 0 527 29 561
rect 63 527 92 561
rect 0 526 92 527
rect 0 17 92 21
rect 0 -17 29 17
rect 63 -17 92 17
<< viali >>
rect 29 527 63 561
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fill_1
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 92 592 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 92 48 1 VGND
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 92 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__fill_1.gds
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 92 214
string MASKHINTS_NSDM 0 -38 92 204
string MASKHINTS_PSDM 0 272 92 582
<< end >>
