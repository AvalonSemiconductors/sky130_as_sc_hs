magic
tech sky130A
magscale 1 2
timestamp 1740589929
<< nwell >>
rect -38 262 1786 582
<< pwell >>
rect 0 34 1748 204
rect 0 24 1104 34
rect 0 22 736 24
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 190 298 220 496
rect 432 298 462 496
rect 528 298 558 496
rect 624 298 654 496
rect 948 298 978 496
rect 1024 298 1054 496
rect 1344 298 1374 496
rect 1430 298 1460 496
rect 1516 298 1546 496
rect 1602 298 1632 496
<< nmoslvt >>
rect 80 48 110 178
rect 190 48 220 178
rect 432 48 462 144
rect 528 48 558 178
rect 720 48 750 178
rect 948 48 978 178
rect 1132 48 1162 178
rect 1344 48 1374 178
rect 1430 48 1460 178
rect 1516 48 1546 178
rect 1602 48 1632 178
<< ndiff >>
rect 27 166 80 178
rect 27 132 35 166
rect 69 132 80 166
rect 27 48 80 132
rect 110 98 190 178
rect 110 64 130 98
rect 164 64 190 98
rect 110 48 190 64
rect 220 166 310 178
rect 220 132 268 166
rect 302 132 310 166
rect 488 144 528 178
rect 220 48 310 132
rect 364 132 432 144
rect 364 98 373 132
rect 407 98 432 132
rect 364 48 432 98
rect 462 98 528 144
rect 462 64 473 98
rect 507 64 528 98
rect 462 48 528 64
rect 558 48 720 178
rect 750 166 840 178
rect 750 132 798 166
rect 832 132 840 166
rect 750 48 840 132
rect 894 98 948 178
rect 894 64 903 98
rect 937 64 948 98
rect 894 48 948 64
rect 978 48 1132 178
rect 1162 166 1236 178
rect 1162 132 1194 166
rect 1228 132 1236 166
rect 1162 48 1236 132
rect 1290 98 1344 178
rect 1290 64 1299 98
rect 1333 64 1344 98
rect 1290 48 1344 64
rect 1374 166 1430 178
rect 1374 132 1385 166
rect 1419 132 1430 166
rect 1374 48 1430 132
rect 1460 170 1516 178
rect 1460 56 1471 170
rect 1505 56 1516 170
rect 1460 48 1516 56
rect 1546 166 1602 178
rect 1546 132 1557 166
rect 1591 132 1602 166
rect 1546 48 1602 132
rect 1632 170 1721 178
rect 1632 56 1643 170
rect 1677 56 1721 170
rect 1632 48 1721 56
<< pdiff >>
rect 27 476 80 496
rect 27 310 35 476
rect 69 310 80 476
rect 27 298 80 310
rect 110 486 190 496
rect 110 384 132 486
rect 166 384 190 486
rect 110 298 190 384
rect 220 476 310 496
rect 220 310 268 476
rect 302 310 310 476
rect 220 298 310 310
rect 364 476 432 496
rect 364 310 373 476
rect 407 310 432 476
rect 364 298 432 310
rect 462 486 528 496
rect 462 384 473 486
rect 507 384 528 486
rect 462 298 528 384
rect 558 298 624 496
rect 654 476 840 496
rect 654 310 798 476
rect 832 310 840 476
rect 654 298 840 310
rect 894 484 948 496
rect 894 382 903 484
rect 937 382 948 484
rect 894 298 948 382
rect 978 298 1024 496
rect 1054 476 1236 496
rect 1054 310 1194 476
rect 1228 310 1236 476
rect 1054 298 1236 310
rect 1290 484 1344 496
rect 1290 310 1299 484
rect 1333 310 1344 484
rect 1290 298 1344 310
rect 1374 476 1430 496
rect 1374 306 1385 476
rect 1419 306 1430 476
rect 1374 298 1430 306
rect 1460 484 1516 496
rect 1460 372 1471 484
rect 1505 372 1516 484
rect 1460 298 1516 372
rect 1546 476 1602 496
rect 1546 306 1557 476
rect 1591 306 1602 476
rect 1546 298 1602 306
rect 1632 488 1720 496
rect 1632 308 1643 488
rect 1677 308 1720 488
rect 1632 298 1720 308
<< ndiffc >>
rect 35 132 69 166
rect 130 64 164 98
rect 268 132 302 166
rect 373 98 407 132
rect 473 64 507 98
rect 798 132 832 166
rect 903 64 937 98
rect 1194 132 1228 166
rect 1299 64 1333 98
rect 1385 132 1419 166
rect 1471 56 1505 170
rect 1557 132 1591 166
rect 1643 56 1677 170
<< pdiffc >>
rect 35 310 69 476
rect 132 384 166 486
rect 268 310 302 476
rect 373 310 407 476
rect 473 384 507 486
rect 798 310 832 476
rect 903 382 937 484
rect 1194 310 1228 476
rect 1299 310 1333 484
rect 1385 306 1419 476
rect 1471 372 1505 484
rect 1557 306 1591 476
rect 1643 308 1677 488
<< poly >>
rect 80 496 110 522
rect 190 496 220 522
rect 432 496 462 522
rect 528 496 558 522
rect 624 496 654 522
rect 948 496 978 522
rect 1024 496 1054 522
rect 1344 496 1374 522
rect 1430 496 1460 522
rect 1516 496 1546 522
rect 1602 496 1632 522
rect 80 266 110 298
rect 190 266 220 298
rect 432 266 462 298
rect 528 266 558 298
rect 624 266 654 298
rect 80 250 148 266
rect 80 216 104 250
rect 138 216 148 250
rect 80 200 148 216
rect 190 250 244 266
rect 190 216 200 250
rect 234 216 244 250
rect 190 200 244 216
rect 432 250 486 266
rect 432 216 442 250
rect 476 216 486 250
rect 80 178 110 200
rect 190 178 220 200
rect 432 198 486 216
rect 528 250 582 266
rect 528 216 538 250
rect 572 216 582 250
rect 528 198 582 216
rect 624 250 678 266
rect 624 216 634 250
rect 668 216 678 250
rect 624 198 678 216
rect 720 250 774 266
rect 720 216 730 250
rect 764 216 774 250
rect 720 198 774 216
rect 816 250 870 268
rect 948 250 978 298
rect 1024 266 1054 298
rect 816 216 826 250
rect 860 216 978 250
rect 816 200 870 216
rect 432 144 462 198
rect 528 178 558 198
rect 720 178 750 198
rect 948 178 978 216
rect 1020 250 1074 266
rect 1020 216 1030 250
rect 1064 216 1074 250
rect 1020 198 1074 216
rect 1116 250 1170 266
rect 1116 216 1126 250
rect 1160 216 1170 250
rect 1116 198 1170 216
rect 1212 250 1266 266
rect 1212 216 1222 250
rect 1256 248 1266 250
rect 1344 252 1374 298
rect 1430 254 1460 298
rect 1516 254 1546 298
rect 1602 254 1632 298
rect 1430 252 1632 254
rect 1344 248 1632 252
rect 1256 218 1632 248
rect 1256 216 1374 218
rect 1212 214 1374 216
rect 1212 198 1266 214
rect 1132 178 1162 198
rect 1344 178 1374 214
rect 1430 178 1460 218
rect 1516 216 1632 218
rect 1516 178 1546 216
rect 1602 178 1632 216
rect 80 22 110 48
rect 190 22 220 48
rect 432 22 462 48
rect 528 22 558 48
rect 720 22 750 48
rect 948 22 978 48
rect 1132 22 1162 48
rect 1344 22 1374 48
rect 1430 22 1460 48
rect 1516 22 1546 48
rect 1602 22 1632 48
<< polycont >>
rect 104 216 138 250
rect 200 216 234 250
rect 442 216 476 250
rect 538 216 572 250
rect 634 216 668 250
rect 730 216 764 250
rect 826 216 860 250
rect 1030 216 1064 250
rect 1126 216 1160 250
rect 1222 216 1256 250
<< locali >>
rect 0 561 1748 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 526 1748 527
rect 35 476 69 492
rect 132 486 166 526
rect 132 368 166 384
rect 268 476 302 492
rect 35 166 69 310
rect 104 250 154 266
rect 138 216 154 250
rect 104 200 154 216
rect 200 250 234 266
rect 200 166 234 216
rect 69 132 200 166
rect 268 166 302 310
rect 35 116 69 132
rect 268 116 302 132
rect 373 476 407 492
rect 473 486 507 526
rect 473 368 507 384
rect 798 476 832 492
rect 373 166 407 310
rect 903 484 937 526
rect 903 366 937 382
rect 1194 476 1228 492
rect 798 268 832 310
rect 442 250 498 266
rect 476 216 498 250
rect 442 200 498 216
rect 538 250 572 266
rect 538 166 572 216
rect 634 250 668 266
rect 634 198 668 216
rect 730 250 764 266
rect 730 198 764 216
rect 798 250 860 268
rect 1194 266 1228 310
rect 1299 484 1333 526
rect 1299 286 1333 310
rect 1385 476 1419 492
rect 1471 484 1505 526
rect 1471 356 1505 372
rect 1557 476 1591 492
rect 1419 306 1484 318
rect 1385 284 1484 306
rect 1557 284 1591 306
rect 1643 488 1677 526
rect 1643 292 1677 308
rect 798 216 826 250
rect 798 200 860 216
rect 1030 250 1064 266
rect 373 132 572 166
rect 798 166 832 200
rect 1030 198 1064 216
rect 1126 250 1160 266
rect 1126 198 1160 216
rect 1194 250 1256 266
rect 1194 216 1222 250
rect 1194 198 1256 216
rect 1385 246 1591 284
rect 1385 220 1484 246
rect 798 116 832 132
rect 1194 166 1228 198
rect 1194 116 1228 132
rect 1385 166 1419 220
rect 1385 116 1419 132
rect 1471 170 1505 186
rect 112 64 130 98
rect 164 64 180 98
rect 373 82 407 98
rect 456 64 473 98
rect 507 64 524 98
rect 886 64 903 98
rect 937 64 954 98
rect 1282 64 1299 98
rect 1333 64 1350 98
rect 130 21 164 64
rect 473 21 507 64
rect 903 21 937 64
rect 1299 21 1333 64
rect 1557 166 1591 246
rect 1557 116 1591 132
rect 1643 170 1677 186
rect 1471 21 1505 56
rect 1643 21 1677 56
rect 0 17 1748 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 268 374 302 408
rect 200 132 234 166
rect 634 216 668 250
rect 730 216 764 250
rect 1030 216 1064 250
rect 1126 216 1160 250
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 256 408 308 416
rect 256 374 268 408
rect 302 374 668 408
rect 256 366 308 374
rect 634 350 668 374
rect 634 316 1160 350
rect 634 266 668 316
rect 1126 266 1160 316
rect 628 250 674 266
rect 628 216 634 250
rect 668 216 674 250
rect 628 204 674 216
rect 724 250 770 262
rect 724 216 730 250
rect 764 216 770 250
rect 724 204 770 216
rect 1020 250 1074 262
rect 1020 216 1030 250
rect 1064 216 1074 250
rect 1020 206 1074 216
rect 1116 250 1170 266
rect 1116 216 1126 250
rect 1160 216 1170 250
rect 194 166 240 178
rect 194 132 200 166
rect 234 132 240 166
rect 194 110 240 132
rect 730 110 764 204
rect 1030 110 1064 206
rect 1116 204 1170 216
rect 194 76 1064 110
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dyn_dfxtp_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1748 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali 119 221 153 255 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel locali 136 238 136 238 0 FreeSans 200 0 0 0 CLK
flabel locali 442 221 476 255 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali 459 238 459 238 0 FreeSans 200 0 0 0 D
flabel locali 1428 221 1462 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali 1445 238 1445 238 0 FreeSans 200 0 0 0 Q
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__dyn_dfxtp_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 1748 220
string MASKHINTS_NSDM 0 -38 1748 209
string MASKHINTS_PSDM 0 273 1748 582
<< end >>
