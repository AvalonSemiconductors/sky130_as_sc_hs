magic
tech sky130A
magscale 1 2
timestamp 1740314482
<< nwell >>
rect -38 262 590 582
<< pwell >>
rect 6 48 544 204
rect 6 42 362 48
rect 22 26 90 42
rect 22 22 110 26
rect 22 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 168 298 198 496
rect 256 298 286 496
rect 344 298 374 496
rect 432 298 462 496
<< nmoslvt >>
rect 80 48 110 178
rect 168 48 198 178
rect 256 48 286 178
rect 344 48 374 178
rect 432 48 462 178
<< ndiff >>
rect 27 140 80 178
rect 27 106 35 140
rect 69 106 80 140
rect 27 48 80 106
rect 110 92 168 178
rect 110 58 121 92
rect 155 58 168 92
rect 110 48 168 58
rect 198 144 256 178
rect 198 110 210 144
rect 244 110 256 144
rect 198 48 256 110
rect 286 170 344 178
rect 286 64 298 170
rect 332 64 344 170
rect 286 48 344 64
rect 374 170 432 178
rect 374 136 386 170
rect 420 136 432 170
rect 374 48 432 136
rect 462 170 522 178
rect 462 57 476 170
rect 510 57 522 170
rect 462 48 522 57
<< pdiff >>
rect 27 466 80 496
rect 27 358 35 466
rect 69 358 80 466
rect 27 298 80 358
rect 110 488 168 496
rect 110 426 121 488
rect 155 426 168 488
rect 110 298 168 426
rect 198 432 256 496
rect 198 398 210 432
rect 244 398 256 432
rect 198 298 256 398
rect 286 488 344 496
rect 286 354 298 488
rect 332 354 344 488
rect 286 298 344 354
rect 374 474 432 496
rect 374 343 386 474
rect 420 343 432 474
rect 374 298 432 343
rect 462 488 520 496
rect 462 354 474 488
rect 508 354 520 488
rect 462 298 520 354
<< ndiffc >>
rect 35 106 69 140
rect 121 58 155 92
rect 210 110 244 144
rect 298 64 332 170
rect 386 136 420 170
rect 476 57 510 170
<< pdiffc >>
rect 35 358 69 466
rect 121 426 155 488
rect 210 398 244 432
rect 298 354 332 488
rect 386 343 420 474
rect 474 354 508 488
<< poly >>
rect 80 496 110 522
rect 168 496 198 522
rect 256 496 286 522
rect 344 496 374 522
rect 432 496 462 522
rect 80 260 110 298
rect 168 266 198 298
rect 28 250 110 260
rect 28 216 44 250
rect 78 216 110 250
rect 28 200 110 216
rect 80 178 110 200
rect 152 256 206 266
rect 256 264 286 298
rect 344 282 374 298
rect 432 282 462 298
rect 344 264 462 282
rect 256 256 462 264
rect 152 250 462 256
rect 152 216 162 250
rect 196 248 462 250
rect 196 232 374 248
rect 196 222 286 232
rect 196 216 206 222
rect 152 198 206 216
rect 168 178 198 198
rect 256 178 286 222
rect 344 178 374 232
rect 432 178 462 248
rect 80 22 110 48
rect 168 22 198 48
rect 256 22 286 48
rect 344 22 374 48
rect 432 22 462 48
<< polycont >>
rect 44 216 78 250
rect 162 216 196 250
<< locali >>
rect 0 561 552 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 526 552 527
rect 121 488 155 526
rect 35 466 69 484
rect 298 488 332 526
rect 121 410 155 426
rect 210 432 264 448
rect 244 398 264 432
rect 210 382 264 398
rect 69 358 176 376
rect 35 342 176 358
rect 31 250 84 296
rect 31 216 44 250
rect 78 216 84 250
rect 31 200 84 216
rect 142 276 176 342
rect 230 304 264 382
rect 298 338 332 354
rect 386 474 420 490
rect 386 304 420 343
rect 474 488 508 526
rect 474 338 508 354
rect 142 250 196 276
rect 142 216 162 250
rect 142 198 196 216
rect 230 242 420 304
rect 142 166 176 198
rect 35 140 176 166
rect 230 160 264 242
rect 69 132 176 140
rect 210 144 264 160
rect 35 90 69 106
rect 244 110 264 144
rect 104 92 172 98
rect 210 94 264 110
rect 298 170 332 188
rect 104 58 121 92
rect 155 58 172 92
rect 386 170 420 242
rect 386 120 420 136
rect 476 170 510 188
rect 121 21 155 58
rect 298 21 332 64
rect 476 21 510 57
rect 0 17 552 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buff_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 552 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 34 255 68 289 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 51 272 51 272 0 FreeSans 200 0 0 0 A
flabel locali s 238 255 272 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 255 272 255 272 0 FreeSans 200 0 0 0 Y
flabel locali 357 255 391 289 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali 374 272 374 272 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__buff_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 552 216
string MASKHINTS_NSDM 0 -38 552 204
string MASKHINTS_PSDM 0 272 552 582
<< end >>
