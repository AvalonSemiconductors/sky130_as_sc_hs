magic
tech sky130A
magscale 1 2
timestamp 1739961801
<< nwell >>
rect -38 262 958 582
<< pwell >>
rect 0 28 920 204
rect 0 22 736 28
rect 26 -20 90 22
<< pmos >>
rect 80 298 110 496
rect 166 298 196 496
rect 260 298 290 496
rect 350 298 380 496
rect 540 298 570 496
rect 626 298 656 496
rect 712 298 742 496
rect 798 298 828 496
<< nmoslvt >>
rect 80 48 110 178
rect 166 48 196 178
rect 260 48 290 178
rect 344 48 374 178
rect 540 48 570 178
rect 626 48 656 178
rect 712 48 742 178
rect 798 48 828 178
<< ndiff >>
rect 27 150 80 178
rect 27 72 35 150
rect 69 72 80 150
rect 27 48 80 72
rect 110 48 166 178
rect 196 92 260 178
rect 196 58 209 92
rect 243 58 260 92
rect 196 48 260 58
rect 290 48 344 178
rect 374 166 433 178
rect 374 76 385 166
rect 419 76 433 166
rect 374 48 433 76
rect 487 150 540 178
rect 487 60 495 150
rect 529 60 540 150
rect 487 48 540 60
rect 570 170 626 178
rect 570 72 581 170
rect 615 72 626 170
rect 570 48 626 72
rect 656 166 712 178
rect 656 60 667 166
rect 701 60 712 166
rect 656 48 712 60
rect 742 170 798 178
rect 742 72 753 170
rect 787 72 798 170
rect 742 48 798 72
rect 828 170 893 178
rect 828 56 841 170
rect 875 56 893 170
rect 828 48 893 56
<< pdiff >>
rect 27 476 80 496
rect 27 422 35 476
rect 69 422 80 476
rect 27 298 80 422
rect 110 488 166 496
rect 110 454 121 488
rect 155 454 166 488
rect 110 298 166 454
rect 196 462 260 496
rect 196 428 209 462
rect 243 428 260 462
rect 196 298 260 428
rect 290 408 350 496
rect 290 374 304 408
rect 338 374 350 408
rect 290 298 350 374
rect 380 476 433 496
rect 380 442 391 476
rect 425 442 433 476
rect 380 298 433 442
rect 487 484 540 496
rect 487 318 495 484
rect 529 318 540 484
rect 487 298 540 318
rect 570 476 626 496
rect 570 306 581 476
rect 615 306 626 476
rect 570 298 626 306
rect 656 484 712 496
rect 656 310 667 484
rect 701 310 712 484
rect 656 298 712 310
rect 742 476 798 496
rect 742 306 753 476
rect 787 306 798 476
rect 742 298 798 306
rect 828 488 893 496
rect 828 306 841 488
rect 875 306 893 488
rect 828 298 893 306
<< ndiffc >>
rect 35 72 69 150
rect 209 58 243 92
rect 385 76 419 166
rect 495 60 529 150
rect 581 72 615 170
rect 667 60 701 166
rect 753 72 787 170
rect 841 56 875 170
<< pdiffc >>
rect 35 422 69 476
rect 121 454 155 488
rect 209 428 243 462
rect 304 374 338 408
rect 391 442 425 476
rect 495 318 529 484
rect 581 306 615 476
rect 667 310 701 484
rect 753 306 787 476
rect 841 306 875 488
<< poly >>
rect 80 496 110 522
rect 166 496 196 522
rect 260 496 290 522
rect 350 496 380 522
rect 540 496 570 522
rect 626 496 656 522
rect 712 496 742 522
rect 798 496 828 522
rect 80 268 110 298
rect 166 268 196 298
rect 260 268 290 298
rect 350 268 380 298
rect 540 268 570 298
rect 42 250 110 268
rect 42 216 52 250
rect 86 216 110 250
rect 42 200 110 216
rect 152 250 206 268
rect 152 216 162 250
rect 196 216 206 250
rect 152 200 206 216
rect 248 250 302 268
rect 248 216 258 250
rect 292 216 302 250
rect 248 200 302 216
rect 344 250 398 268
rect 344 216 354 250
rect 388 216 398 250
rect 344 200 398 216
rect 458 250 570 268
rect 458 216 472 250
rect 506 236 570 250
rect 626 236 656 298
rect 712 236 742 298
rect 798 236 828 298
rect 506 216 828 236
rect 458 200 828 216
rect 80 178 110 200
rect 166 178 196 200
rect 260 178 290 200
rect 344 178 374 200
rect 540 178 570 200
rect 626 178 656 200
rect 712 178 742 200
rect 798 178 828 200
rect 80 22 110 48
rect 166 22 196 48
rect 260 22 290 48
rect 344 22 374 48
rect 540 22 570 48
rect 626 22 656 48
rect 712 22 742 48
rect 798 22 828 48
<< polycont >>
rect 52 216 86 250
rect 162 216 196 250
rect 258 216 292 250
rect 354 216 388 250
rect 472 216 506 250
<< locali >>
rect 0 561 920 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 526 920 527
rect 35 476 69 492
rect 121 488 155 526
rect 104 454 121 488
rect 155 454 172 488
rect 209 476 425 492
rect 209 462 391 476
rect 35 420 69 422
rect 243 458 391 462
rect 209 420 243 428
rect 391 426 425 442
rect 495 484 529 526
rect 35 386 243 420
rect 304 408 338 424
rect 304 366 338 374
rect 42 268 86 352
rect 152 268 198 352
rect 232 268 270 352
rect 304 332 456 366
rect 422 268 456 332
rect 495 302 529 318
rect 581 476 615 492
rect 581 298 615 306
rect 667 484 701 526
rect 42 250 96 268
rect 42 216 52 250
rect 86 216 96 250
rect 42 200 96 216
rect 152 250 196 268
rect 152 216 162 250
rect 232 250 292 268
rect 232 238 258 250
rect 152 200 196 216
rect 248 216 258 238
rect 248 200 292 216
rect 328 250 388 268
rect 328 216 354 250
rect 328 200 388 216
rect 422 250 506 268
rect 422 216 472 250
rect 422 200 506 216
rect 564 254 622 298
rect 667 288 701 310
rect 753 476 787 492
rect 753 254 787 306
rect 841 488 875 526
rect 841 288 875 306
rect 564 220 787 254
rect 422 166 456 200
rect 564 184 622 220
rect 581 170 615 184
rect 35 150 385 166
rect 69 132 385 150
rect 35 56 69 72
rect 192 92 260 96
rect 192 58 209 92
rect 243 58 260 92
rect 419 132 456 166
rect 495 150 529 166
rect 385 60 419 76
rect 209 21 243 58
rect 495 21 529 60
rect 581 56 615 72
rect 667 166 701 186
rect 667 21 701 60
rect 753 170 787 220
rect 753 56 787 72
rect 841 170 875 186
rect 841 21 875 56
rect 0 17 920 21
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ao22_4
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 3 nsew power bidirectional abutment
flabel locali s 51 204 85 238 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 68 221 68 221 0 FreeSans 200 0 0 0 A
flabel locali s 255 204 289 238 0 FreeSans 200 0 0 0 C
port 6 nsew signal input
flabel locali s 272 221 272 221 0 FreeSans 200 0 0 0 C
flabel locali s 153 204 187 238 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel locali s 170 221 170 221 0 FreeSans 200 0 0 0 B
flabel locali s 340 204 374 238 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel locali s 357 221 357 221 0 FreeSans 200 0 0 0 D
flabel locali s 578 204 612 238 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 595 221 595 221 0 FreeSans 200 0 0 0 Y
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_as_sc_hs/gds/sky130_as_sc_hs__ao22_4.gds
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string MASKHINTS_LVTN 0 -4 920 220
string MASKHINTS_NSDM 0 -38 920 209
string MASKHINTS_PSDM 0 273 920 582
<< end >>
