magic
tech sky130A
magscale 1 2
timestamp 1732639285
<< nwell >>
rect -38 262 406 582
<< pwell >>
rect 22 48 346 204
rect 26 44 320 48
rect 26 -20 90 44
<< locali >>
rect 0 526 8 562
rect 360 526 368 562
rect 0 -15 8 21
rect 360 -15 368 21
<< viali >>
rect 8 526 360 562
rect 8 -15 360 21
<< metal1 >>
rect 0 562 368 592
rect 0 526 8 562
rect 360 526 368 562
rect 0 496 368 526
rect 0 21 368 48
rect 0 -15 8 21
rect 360 -15 368 21
rect 0 -48 368 -15
<< labels >>
rlabel comment s 0 0 0 0 4 aaaaaaa
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 1 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 0 -48 368 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 0 496 368 592 1 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
